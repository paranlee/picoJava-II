/****************************************************************
 ---------------------------------------------------------------
     Copyright 1999 Sun Microsystems, Inc., 901 San Antonio
     Road, Palo Alto, CA 94303, U.S.A.  All Rights Reserved.
     The contents of this file are subject to the current
     version of the Sun Community Source License, picoJava-II
     Core ("the License").  You may not use this file except
     in compliance with the License.  You may obtain a copy
     of the License by searching for "Sun Community Source
     License" on the World Wide Web at http://www.sun.com.
     See the License for the rights, obligations, and
     limitations governing use of the contents of this file.

     Sun, Sun Microsystems, the Sun logo, and all Sun-based
     trademarks and logos, Java, picoJava, and all Java-based
     trademarks and logos are trademarks or registered trademarks 
     of Sun Microsystems, Inc. in the United States and other
     countries.
 ----------------------------------------------------------------
******************************************************************/

/* ********************************************************************
 * The ibuf_monitor module monitors icu_vld_d (valid byte),  
 * iu_shift_d (# of read byte), and ic_fill_sel[15:0], 
 * and performs the following tasks:
 *
 * 1) Monitor the ibuffer state at each cycle.   
 * 2) Set flag for each ibuffer state(pattern).
 * 3) Any pattern that does not match the specified group of
 *    patterns will flag an Error and stop the simulation.   
 * 
 * Note: 
 *       1. If the occurrence of a pattern is "0" then the designer
 *          needs to write a specific test to produce the pattern 
 *          so the coverage for ibuf verification can reach 100%.
 *
 *       2. If a specific pattern produced does not fall under
 *          the group, the simulation will be stopped. The designer
 *          must debug it!  
 *	      
 *       3. Boot Mode is not tested by this monitor.
 *
 * Included below is the group of all states(patterns) the ibuffer 
 * may present according to the specs.:
 * 
 * 
 *  	# of valid byte		# of read bytes     Write from Nth byte
 *  	valid[15:0]   		iu_shift_d[7:0]     ic_fill_sel[15:0]
 *
 * Pattern
 * _name:
 *
 * v0r0w0:0000000000000000  (0)	 00000001  (0)	    1111111111111111  (0)
 * v1r0w1:0000000000000001  (1)  00000001  (0)      1111111111111110  (1)
 * v1r1w0:0000000000000001  (1)  00000010  (1)      1111111111111111  (0)
 * v2r0w2:0000000000000011  (2)  00000001  (0)      1111111111111100  (2)
 * v2r1w1:0000000000000011  (2)  00000010  (1)      1111111111111110  (1)
 * v2r2w0:0000000000000011  (2)  00000100  (2)      1111111111111111  (0)
 * v3r0w3:0000000000000111  (3)  00000001  (0)      1111111111111000  (3)
 * v3r1w2:0000000000000111  (3)  00000010  (1)      1111111111111100  (2)
 * v3r2w1:0000000000000111  (3)  00000100  (2)      1111111111111110  (1)
 * v3r3w0:0000000000000111  (3)  00001000  (3)      1111111111111111  (0)
 * v4r0w4:0000000000001111  (4)  00000001  (0)      1111111111110000  (4)
 * v4r1w3:0000000000001111  (4)  00000010  (1)      1111111111111000  (3)
 * v4r2w2:0000000000001111  (4)  00000100  (2)      1111111111111100  (2)
 * v4r3w1:0000000000001111  (4)  00001000  (3)      1111111111111110  (1)
 * v4r4w0:0000000000001111  (4)  00010000  (4)      1111111111111111  (0)
 * v5r0w5:0000000000011111  (5)  00000001  (0)      1111111111100000  (5)
 * v5r1w4:0000000000011111  (5)  00000010  (1)      1111111111110000  (4)
 * v5r2w3:0000000000011111  (5)  00000100  (2)      1111111111111000  (3)
 * v5r3w2:0000000000011111  (5)  00001000  (3)      1111111111111100  (2)
 * v5r4w1:0000000000011111  (5)  00010000  (4)      1111111111111110  (1)
 * v5r5w0:0000000000011111  (5)  00100000  (5)      1111111111111111  (0)
 * v6r0w6:0000000000111111  (6)  00000001  (0)      1111111111000000  (6)
 * v6r1w5:0000000000111111  (6)  00000010  (1)      1111111111100000  (5)
 * v6r2w4:0000000000111111  (6)  00000100  (2)      1111111111110000  (4)
 * v6r3w3:0000000000111111  (6)  00001000  (3)      1111111111111000  (3)
 * v6r4w2:0000000000111111  (6)  00010000  (4)      1111111111111100  (2)
 * v6r5w1:0000000000111111  (6)  00100000  (5)      1111111111111110  (1)
 **v6r6w0:0000000000111111  (6)  01000000  (6)      1111111111111111  (0)
 * v7r0w7:0000000001111111  (7)  00000001  (0)      1111111110000000  (7)
 * v7r1w6:0000000001111111  (7)  00000010  (1)      1111111111000000  (6)
 * v7r2w5:0000000001111111  (7)  00000100  (2)      1111111111100000  (5)
 * v7r3w4:0000000001111111  (7)  00001000  (3)      1111111111110000  (4)
 * v7r4w3:0000000001111111  (7)  00010000  (4)      1111111111111000  (3)
 * v7r5w2:0000000001111111  (7)  00100000  (5)      1111111111111100  (2)
 **v7r6w1:0000000001111111  (7)  01000000  (6)      1111111111111110  (1)
 **v7r7w0:0000000001111111  (7)  10000000  (7)      1111111111111111  (0)
 * v8r0w8:0000000011111111  (8)  00000001  (0)      1111111100000000  (8)
 * v8r1w7:0000000011111111  (8)  00000010  (1)      1111111110000000  (7)
 * v8r2w6:0000000011111111  (8)  00000100  (2)      1111111111000000  (6)
 * v8r3w5:0000000011111111  (8)  00001000  (3)      1111111111100000  (5)
 * v8r4w4:0000000011111111  (8)  00010000  (4)      1111111111110000  (4)
 * v8r5w3:0000000011111111  (8)  00100000  (5)      1111111111111000  (3)
 **v8r6w2:0000000011111111  (8)  01000000  (6)      1111111111111100  (2)
 **v8r7w1:0000000011111111  (8)  10000000  (7)      1111111111111110  (1)
 * v9r0w9:0000000111111111  (9)  00000001  (0)      1111111000000000  (9)
 * v9r1w8:0000000111111111  (9)  00000010  (1)      1111111100000000  (8)
 * v9r2w7:0000000111111111  (9)  00000100  (2)      1111111110000000  (7)
 * v9r3w6:0000000111111111  (9)  00001000  (3)      1111111111000000  (6)
 * v9r4w5:0000000111111111  (9)  00010000  (4)      1111111111100000  (5)
 * v9r5w4:0000000111111111  (9)  00100000  (5)      1111111111110000  (4)
 **v9r6w3:0000000111111111  (9)  01000000  (6)      1111111111111000  (3)
 **v9r7w2:0000000111111111  (9)  10000000  (7)      1111111111111100  (2)
 * vAr0wA:0000001111111111  (A)  00000001  (0)      1111110000000000  (A)
 * vAr1w9:0000001111111111  (A)  00000010  (1)      1111111000000000  (9)
 * vAr2w8:0000001111111111  (A)  00000100  (2)      1111111100000000  (8)
 * vAr3w7:0000001111111111  (A)  00001000  (3)      1111111110000000  (7)
 * vAr4w6:0000001111111111  (A)  00010000  (4)      1111111111000000  (6)
 * vAr5w5:0000001111111111  (A)  00100000  (5)      1111111111100000  (5)
 **vAr6w4:0000001111111111  (A)  01000000  (6)      1111111111110000  (4)
 **vAr7w3:0000001111111111  (A)  10000000  (7)      1111111111111000  (3)
 * vBr0wB:0000011111111111  (B)  00000001  (0)      1111100000000000  (B)
 * vBr1wA:0000011111111111  (B)  00000010  (1)      1111110000000000  (A)
 * vBr2w9:0000011111111111  (B)  00000100  (2)      1111111000000000  (9)
 * vBr3w8:0000011111111111  (B)  00001000  (3)      1111111100000000  (8)
 * vBr4w7:0000011111111111  (B)  00010000  (4)      1111111110000000  (7)
 * vBr5w6:0000011111111111  (B)  00100000  (5)      1111111111000000  (6)
 **vBr6w5:0000011111111111  (B)  01000000  (6)      1111111111100000  (5)
 **vBr7w4:0000011111111111  (B)  10000000  (7)      1111111111110000  (4)
 * vCr0wC:0000111111111111  (C)  00000001  (0)      1111000000000000  (C)
 * vCr1wB:0000111111111111  (C)  00000010  (1)      1111100000000000  (B)
 * vCr2wA:0000111111111111  (C)  00000100  (2)      1111110000000000  (A)
 * vCr3w9:0000111111111111  (C)  00001000  (3)      1111111000000000  (9)
 * vCr4w8:0000111111111111  (C)  00010000  (4)      1111111100000000  (8)
 * vCr5w7:0000111111111111  (C)  00100000  (5)      1111111110000000  (7)
 **vCr6w6:0000111111111111  (C)  01000000  (6)      1111111111000000  (6)
 **vCr7w5:0000111111111111  (C)  10000000  (7)      1111111111100000  (5)
 **vDr0wD:0001111111111111  (D)  00000001  (0)      1110000000000000  (D)
 **vDr1wC:0001111111111111  (D)  00000010  (1)      1111000000000000  (C)
 **vDr2wB:0001111111111111  (D)  00000100  (2)      1111100000000000  (B)
 **vDr3wA:0001111111111111  (D)  00001000  (3)      1111110000000000  (A)
 **vDr4w9:0001111111111111  (D)  00010000  (4)      1111111000000000  (9)
 **vDr5w8:0001111111111111  (D)  00100000  (5)      1111111100000000  (8)
 **vDr6w7:0001111111111111  (D)  01000000  (6)      1111111110000000  (7)
 **vDr7w6:0001111111111111  (D)  10000000  (7)      1111111111000000  (6)
 **vEr0wE:0011111111111111  (E)  00000001  (0)      1100000000000000  (E)
 **vEr1wD:0011111111111111  (E)  00000010  (1)      1110000000000000  (D)
 **vEr2wC:0011111111111111  (E)  00000100  (2)      1111000000000000  (C)
 **vEr3wB:0011111111111111  (E)  00001000  (3)      1111100000000000  (B)
 **vEr4wA:0011111111111111  (E)  00010000  (4)      1111110000000000  (A)
 **vEr5w9:0011111111111111  (E)  00100000  (5)      1111111000000000  (9)
 **vEr6w8:0011111111111111  (E)  01000000  (6)      1111111100000000  (8)
 **vEr7w7:0011111111111111  (E)  10000000  (7)      1111111110000000  (7)
 **vFr0wF:0111111111111111  (F)  00000001  (0)      1000000000000000  (F)
 **vFr1wE:0111111111111111  (F)  00000010  (1)      1100000000000000  (E)
 **vFr2wD:0111111111111111  (F)  00000100  (2)      1110000000000000  (D)
 **vFr3wC:0111111111111111  (F)  00001000  (3)      1111000000000000  (C)
 **vFr4wB:0111111111111111  (F)  00010000  (4)      1111100000000000  (B)
 **vFr5wA:0111111111111111  (F)  00100000  (5)      1111110000000000  (A)
 **vFr6w9:0111111111111111  (F)  01000000  (6)      1111111000000000  (9)
 **vFr7w8:0111111111111111  (F)  10000000  (7)      1111111100000000  (8)
 **vGr0wG:1111111111111111  (G)  00000001  (0)      0000000000000000  (G)
 **vGr1wF:1111111111111111  (G)  00000010  (1)      1000000000000000  (F)
 **vGr2wE:1111111111111111  (G)  00000100  (2)      1100000000000000  (E)
 **vGr3wD:1111111111111111  (G)  00001000  (3)      1110000000000000  (D)
 **vGr4wC:1111111111111111  (G)  00010000  (4)      1111000000000000  (C)
 **vGr5wB:1111111111111111  (G)  00100000  (5)      1111100000000000  (B)
 **vGr6wA:1111111111111111  (G)  01000000  (6)      1111110000000000  (A)
 **vGr7w9:1111111111111111  (G)  10000000  (7)      1111111000000000  (9)
 *
 * ***************************************************************** */

module ibuf_monitor(
        clk,
        num_val_byte,
        num_rd_byte,
        nth_wr_byte_input,
        reset
	);

input		clk, reset;	
input  	[15:0]	num_val_byte;	
input  	[7:0]	num_rd_byte;	
input  	[15:0]	nth_wr_byte_input;	

reg	[15:0]	nth_wr_byte;
always @(nth_wr_byte_input or num_rd_byte or num_val_byte) begin
  case(num_rd_byte)
    8'b00000001: nth_wr_byte = nth_wr_byte_input;
    8'b00000010: nth_wr_byte = (nth_wr_byte_input >> 1) | 32'h8000;
    8'b00000100: nth_wr_byte = (nth_wr_byte_input >> 2) | 32'hc000;
    8'b00001000: nth_wr_byte = (nth_wr_byte_input >> 3) | 32'he000;
    8'b00010000: nth_wr_byte = (nth_wr_byte_input >> 4) | 32'hf000;
    8'b00100000: nth_wr_byte = (nth_wr_byte_input >> 5) | 32'hf800;
    8'b01000000: nth_wr_byte = (nth_wr_byte_input >> 6) | 32'hfc00;
    8'b10000000: nth_wr_byte = (nth_wr_byte_input >> 7) | 32'hfe00;
  endcase
end

reg
  v0r0w0, v1r0w1, v1r1w0, v2r0w2, v2r1w1, v2r2w0, v3r0w3, v3r1w2,
  v3r2w1, v3r3w0, v4r0w4, v4r1w3, v4r2w2, v4r3w1, v4r4w0, v5r0w5,
  v5r1w4, v5r2w3, v5r3w2, v5r4w1, v5r5w0, v6r0w6, v6r1w5, v6r2w4,
  v6r3w3, v6r4w2, v6r5w1, v6r6w0, v7r0w7, v7r1w6, v7r2w5, v7r3w4,
  v7r4w3, v7r5w2, v7r6w1, v7r7w0, v8r0w8, v8r1w7, v8r2w6, v8r3w5,
  v8r4w4, v8r5w3, v8r6w2, v8r7w1, v9r0w9, v9r1w8, v9r2w7, v9r3w6,
  v9r4w5, v9r5w4, v9r6w3, v9r7w2, vAr0wA, vAr1w9, vAr2w8, vAr3w7,
  vAr4w6, vAr5w5, vAr6w4, vAr7w3, vBr0wB, vBr1wA, vBr2w9, vBr3w8,
  vBr4w7, vBr5w6, vBr6w5, vBr7w4, vCr0wC, vCr1wB, vCr2wA, vCr3w9,
  vCr4w8, vCr5w7, vCr6w6, vCr7w5, vDr0wD, vDr1wC, vDr2wB, vDr3wA,
  vDr4w9, vDr5w8, vDr6w7, vDr7w6, vEr0wE, vEr1wD, vEr2wC, vEr3wB,
  vEr4wA, vEr5w9, vEr6w8, vEr7w7, vFr0wF, vFr1wE, vFr2wD, vFr3wC,
  vFr4wB, vFr5wA, vFr6w9, vFr7w8, vGr0wG, vGr1wF, vGr2wE, vGr3wD,
  vGr4wC, vGr5wB, vGr6wA, vGr7w9;


wire 	[39:0]  ibuf_pattern = {num_val_byte,num_rd_byte,nth_wr_byte}; 

integer mcd;
integer monitor_enable;

initial begin

  v0r0w0 = 0; v1r0w1 = 0; v1r1w0 = 0; v2r0w2 = 0; v2r1w1 = 0;
  v2r2w0 = 0; v3r0w3 = 0; v3r1w2 = 0; v3r2w1 = 0; v3r3w0 = 0;
  v4r0w4 = 0; v4r1w3 = 0; v4r2w2 = 0; v4r3w1 = 0; v4r4w0 = 0;
  v5r0w5 = 0; v5r1w4 = 0; v5r2w3 = 0; v5r3w2 = 0; v5r4w1 = 0;
  v5r5w0 = 0; v6r0w6 = 0; v6r1w5 = 0; v6r2w4 = 0; v6r3w3 = 0;
  v6r4w2 = 0; v6r5w1 = 0; v6r6w0 = 0; v7r0w7 = 0; v7r1w6 = 0;
  v7r2w5 = 0; v7r3w4 = 0; v7r4w3 = 0; v7r5w2 = 0; v7r6w1 = 0;
  v7r7w0 = 0; v8r0w8 = 0; v8r1w7 = 0; v8r2w6 = 0; v8r3w5 = 0;
  v8r4w4 = 0; v8r5w3 = 0; v8r6w2 = 0; v8r7w1 = 0; v9r0w9 = 0;
  v9r1w8 = 0; v9r2w7 = 0; v9r3w6 = 0; v9r4w5 = 0; v9r5w4 = 0;
  v9r6w3 = 0; v9r7w2 = 0; vAr0wA = 0; vAr1w9 = 0; vAr2w8 = 0;
  vAr3w7 = 0; vAr4w6 = 0; vAr5w5 = 0; vAr6w4 = 0; vAr7w3 = 0;
  vBr0wB = 0; vBr1wA = 0; vBr2w9 = 0; vBr3w8 = 0; vBr4w7 = 0;
  vBr5w6 = 0; vBr6w5 = 0; vBr7w4 = 0; vCr0wC = 0; vCr1wB = 0;
  vCr2wA = 0; vCr3w9 = 0; vCr4w8 = 0; vCr5w7 = 0; vCr6w6 = 0;
  vCr7w5 = 0; vDr0wD = 0; vDr1wC = 0; vDr2wB = 0; vDr3wA = 0;
  vDr4w9 = 0; vDr5w8 = 0; vDr6w7 = 0; vDr7w6 = 0; vEr0wE = 0;
  vEr1wD = 0; vEr2wC = 0; vEr3wB = 0; vEr4wA = 0; vEr5w9 = 0;
  vEr6w8 = 0; vEr7w7 = 0; vFr0wF = 0; vFr1wE = 0; vFr2wD = 0;
  vFr3wC = 0; vFr4wB = 0; vFr5wA = 0; vFr6w9 = 0; vFr7w8 = 0;
  vGr0wG = 0; vGr1wF = 0; vGr2wE = 0; vGr3wD = 0; vGr4wC = 0;
  vGr5wB = 0; vGr6wA = 0; vGr7w9 = 0;

  monitor_enable = ($test$plusargs("ibuf_mon")) ? 1 : 0;

  if (monitor_enable)
    mcd = $fopen("ibuf.dat");

end

always @ (posedge clk)  begin
  if (monitor_enable) begin
    case(ibuf_pattern)
      40'b0000000000000000000000011111111111111111: v0r0w0 = 1'b1;
      40'b0000000000000001000000011111111111111110: v1r0w1 = 1'b1;
      40'b0000000000000001000000101111111111111111: v1r1w0 = 1'b1;
      40'b0000000000000011000000011111111111111100: v2r0w2 = 1'b1;
      40'b0000000000000011000000101111111111111110: v2r1w1 = 1'b1;
      40'b0000000000000011000001001111111111111111: v2r2w0 = 1'b1;
      40'b0000000000000111000000011111111111111000: v3r0w3 = 1'b1;
      40'b0000000000000111000000101111111111111100: v3r1w2 = 1'b1;
      40'b0000000000000111000001001111111111111110: v3r2w1 = 1'b1;
      40'b0000000000000111000010001111111111111111: v3r3w0 = 1'b1;
      40'b0000000000001111000000011111111111110000: v4r0w4 = 1'b1;
      40'b0000000000001111000000101111111111111000: v4r1w3 = 1'b1;
      40'b0000000000001111000001001111111111111100: v4r2w2 = 1'b1;
      40'b0000000000001111000010001111111111111110: v4r3w1 = 1'b1;
      40'b0000000000001111000100001111111111111111: v4r4w0 = 1'b1;
      40'b0000000000011111000000011111111111100000: v5r0w5 = 1'b1;
      40'b0000000000011111000000101111111111110000: v5r1w4 = 1'b1;
      40'b0000000000011111000001001111111111111000: v5r2w3 = 1'b1;
      40'b0000000000011111000010001111111111111100: v5r3w2 = 1'b1;
      40'b0000000000011111000100001111111111111110: v5r4w1 = 1'b1;
      40'b0000000000011111001000001111111111111111: v5r5w0 = 1'b1;
      40'b0000000000111111000000011111111111000000: v6r0w6 = 1'b1;
      40'b0000000000111111000000101111111111100000: v6r1w5 = 1'b1;
      40'b0000000000111111000001001111111111110000: v6r2w4 = 1'b1;
      40'b0000000000111111000010001111111111111000: v6r3w3 = 1'b1;
      40'b0000000000111111000100001111111111111100: v6r4w2 = 1'b1;
      40'b0000000000111111001000001111111111111110: v6r5w1 = 1'b1;
      40'b0000000000111111010000001111111111111111: v6r6w0 = 1'b1;
      40'b0000000001111111000000011111111110000000: v7r0w7 = 1'b1;
      40'b0000000001111111000000101111111111000000: v7r1w6 = 1'b1;
      40'b0000000001111111000001001111111111100000: v7r2w5 = 1'b1;
      40'b0000000001111111000010001111111111110000: v7r3w4 = 1'b1;
      40'b0000000001111111000100001111111111111000: v7r4w3 = 1'b1;
      40'b0000000001111111001000001111111111111100: v7r5w2 = 1'b1;
      40'b0000000001111111010000001111111111111110: v7r6w1 = 1'b1;
      40'b0000000001111111100000001111111111111111: v7r7w0 = 1'b1;
      40'b0000000011111111000000011111111100000000: v8r0w8 = 1'b1;
      40'b0000000011111111000000101111111110000000: v8r1w7 = 1'b1;
      40'b0000000011111111000001001111111111000000: v8r2w6 = 1'b1;
      40'b0000000011111111000010001111111111100000: v8r3w5 = 1'b1;
      40'b0000000011111111000100001111111111110000: v8r4w4 = 1'b1;
      40'b0000000011111111001000001111111111111000: v8r5w3 = 1'b1;
      40'b0000000011111111010000001111111111111100: v8r6w2 = 1'b1;
      40'b0000000011111111100000001111111111111110: v8r7w1 = 1'b1;
      40'b0000000111111111000000011111111000000000: v9r0w9 = 1'b1;
      40'b0000000111111111000000101111111100000000: v9r1w8 = 1'b1;
      40'b0000000111111111000001001111111110000000: v9r2w7 = 1'b1;
      40'b0000000111111111000010001111111111000000: v9r3w6 = 1'b1;
      40'b0000000111111111000100001111111111100000: v9r4w5 = 1'b1;
      40'b0000000111111111001000001111111111110000: v9r5w4 = 1'b1;
      40'b0000000111111111010000001111111111111000: v9r6w3 = 1'b1;
      40'b0000000111111111100000001111111111111100: v9r7w2 = 1'b1;
      40'b0000001111111111000000011111110000000000: vAr0wA = 1'b1;
      40'b0000001111111111000000101111111000000000: vAr1w9 = 1'b1;
      40'b0000001111111111000001001111111100000000: vAr2w8 = 1'b1;
      40'b0000001111111111000010001111111110000000: vAr3w7 = 1'b1;
      40'b0000001111111111000100001111111111000000: vAr4w6 = 1'b1;
      40'b0000001111111111001000001111111111100000: vAr5w5 = 1'b1;
      40'b0000001111111111010000001111111111110000: vAr6w4 = 1'b1;
      40'b0000001111111111100000001111111111111000: vAr7w3 = 1'b1;
      40'b0000011111111111000000011111100000000000: vBr0wB = 1'b1;
      40'b0000011111111111000000101111110000000000: vBr1wA = 1'b1;
      40'b0000011111111111000001001111111000000000: vBr2w9 = 1'b1;
      40'b0000011111111111000010001111111100000000: vBr3w8 = 1'b1;
      40'b0000011111111111000100001111111110000000: vBr4w7 = 1'b1;
      40'b0000011111111111001000001111111111000000: vBr5w6 = 1'b1;
      40'b0000011111111111010000001111111111100000: vBr6w5 = 1'b1;
      40'b0000011111111111100000001111111111110000: vBr7w4 = 1'b1;
      40'b0000111111111111000000011111000000000000: vCr0wC = 1'b1;
      40'b0000111111111111000000101111100000000000: vCr1wB = 1'b1;
      40'b0000111111111111000001001111110000000000: vCr2wA = 1'b1;
      40'b0000111111111111000010001111111000000000: vCr3w9 = 1'b1;
      40'b0000111111111111000100001111111100000000: vCr4w8 = 1'b1;
      40'b0000111111111111001000001111111110000000: vCr5w7 = 1'b1;
      40'b0000111111111111010000001111111111000000: vCr6w6 = 1'b1;
      40'b0000111111111111100000001111111111100000: vCr7w5 = 1'b1;
      40'b0001111111111111000000011110000000000000: vDr0wD = 1'b1;
      40'b0001111111111111000000101111000000000000: vDr1wC = 1'b1;
      40'b0001111111111111000001001111100000000000: vDr2wB = 1'b1;
      40'b0001111111111111000010001111110000000000: vDr3wA = 1'b1;
      40'b0001111111111111000100001111111000000000: vDr4w9 = 1'b1;
      40'b0001111111111111001000001111111100000000: vDr5w8 = 1'b1;
      40'b0001111111111111010000001111111110000000: vDr6w7 = 1'b1;
      40'b0001111111111111100000001111111111000000: vDr7w6 = 1'b1;
      40'b0011111111111111000000011100000000000000: vEr0wE = 1'b1;
      40'b0011111111111111000000101110000000000000: vEr1wD = 1'b1;
      40'b0011111111111111000001001111000000000000: vEr2wC = 1'b1;
      40'b0011111111111111000010001111100000000000: vEr3wB = 1'b1;
      40'b0011111111111111000100001111110000000000: vEr4wA = 1'b1;
      40'b0011111111111111001000001111111000000000: vEr5w9 = 1'b1;
      40'b0011111111111111010000001111111100000000: vEr6w8 = 1'b1;
      40'b0011111111111111100000001111111110000000: vEr7w7 = 1'b1;
      40'b0111111111111111000000011000000000000000: vFr0wF = 1'b1;
      40'b0111111111111111000000101100000000000000: vFr1wE = 1'b1;
      40'b0111111111111111000001001110000000000000: vFr2wD = 1'b1;
      40'b0111111111111111000010001111000000000000: vFr3wC = 1'b1;
      40'b0111111111111111000100001111100000000000: vFr4wB = 1'b1;
      40'b0111111111111111001000001111110000000000: vFr5wA = 1'b1;
      40'b0111111111111111010000001111111000000000: vFr6w9 = 1'b1;
      40'b0111111111111111100000001111111100000000: vFr7w8 = 1'b1;
      40'b1111111111111111000000010000000000000000: vGr0wG = 1'b1;
      40'b1111111111111111000000101000000000000000: vGr1wF = 1'b1;
      40'b1111111111111111000001001100000000000000: vGr2wE = 1'b1;
      40'b1111111111111111000010001110000000000000: vGr3wD = 1'b1;
      40'b1111111111111111000100001111000000000000: vGr4wC = 1'b1;
      40'b1111111111111111001000001111100000000000: vGr5wB = 1'b1;
      40'b1111111111111111010000001111110000000000: vGr6wA = 1'b1;
      40'b1111111111111111100000001111111000000000: vGr7w9 = 1'b1;
      default:
	if (!reset) begin 
	  $display("ERROR: Incorrect ibuf state:");
	  $display("# of valid bytes = %h ;", num_val_byte);
	  $display("# of read  bytes = %h ;", num_rd_byte);
	  $display("Write from Nth byte = %h",nth_wr_byte);
	  $display("Write from Nth byte input = %h", nth_wr_byte_input);
	  $display("*** You must debug this case. ***");
	  $finish;
	end
    endcase
  end
end

always @(`PICOJAVAII.end_of_simulation)
  if(`PICOJAVAII.end_of_simulation & monitor_enable) begin
    $fdisplay(mcd,"vvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvvv");
    $fdisplay(mcd,"0112223333444445555556666666777777778888888899999999AAAAAAAABBBBBBBBCCCCCCCCDDDDDDDDEEEEEEEEFFFFFFFFGGGGGGGG");
    $fdisplay(mcd,"rrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrrr");
    $fdisplay(mcd,"001012012301234012345012345601234567012345670123456701234567012345670123456701234567012345670123456701234567");
    $fdisplay(mcd,"wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww");
    $fdisplay(mcd,"0102103210432105432106543210765432108765432198765432A9876543BA987654CBA98765DCBA9876EDCBA987FEDCBA98GFEDCBA9");
    $fdisplay(mcd," ");
    $fdisplay(mcd,"%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b",
      v0r0w0, v1r0w1, v1r1w0, v2r0w2, v2r1w1, v2r2w0, v3r0w3,
      v3r1w2, v3r2w1, v3r3w0, v4r0w4, v4r1w3, v4r2w2, v4r3w1,
      v4r4w0, v5r0w5, v5r1w4, v5r2w3, v5r3w2, v5r4w1, v5r5w0,
      v6r0w6, v6r1w5, v6r2w4, v6r3w3, v6r4w2, v6r5w1, v6r6w0,
      v7r0w7, v7r1w6, v7r2w5, v7r3w4, v7r4w3, v7r5w2, v7r6w1,
      v7r7w0, v8r0w8, v8r1w7, v8r2w6, v8r3w5, v8r4w4, v8r5w3,
      v8r6w2, v8r7w1, v9r0w9, v9r1w8, v9r2w7, v9r3w6, v9r4w5,
      v9r5w4, v9r6w3, v9r7w2, vAr0wA, vAr1w9, vAr2w8, vAr3w7,
      vAr4w6, vAr5w5, vAr6w4, vAr7w3, vBr0wB, vBr1wA, vBr2w9,
      vBr3w8, vBr4w7, vBr5w6, vBr6w5, vBr7w4, vCr0wC, vCr1wB,
      vCr2wA, vCr3w9, vCr4w8, vCr5w7, vCr6w6, vCr7w5, vDr0wD,
      vDr1wC, vDr2wB, vDr3wA, vDr4w9, vDr5w8, vDr6w7, vDr7w6,
      vEr0wE, vEr1wD, vEr2wC, vEr3wB, vEr4wA, vEr5w9, vEr6w8,
      vEr7w7, vFr0wF, vFr1wE, vFr2wD, vFr3wC, vFr4wB, vFr5wA,
      vFr6w9, vFr7w8, vGr0wG, vGr1wF, vGr2wE, vGr3wD, vGr4wC,
      vGr5wB, vGr6wA, vGr7w9 );
    $display("COVERAGE: ibuffer %b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b",
      v0r0w0, v1r0w1, v1r1w0, v2r0w2, v2r1w1, v2r2w0, v3r0w3,
      v3r1w2, v3r2w1, v3r3w0, v4r0w4, v4r1w3, v4r2w2, v4r3w1,
      v4r4w0, v5r0w5, v5r1w4, v5r2w3, v5r3w2, v5r4w1, v5r5w0,
      v6r0w6, v6r1w5, v6r2w4, v6r3w3, v6r4w2, v6r5w1, v6r6w0,
      v7r0w7, v7r1w6, v7r2w5, v7r3w4, v7r4w3, v7r5w2, v7r6w1,
      v7r7w0, v8r0w8, v8r1w7, v8r2w6, v8r3w5, v8r4w4, v8r5w3,
      v8r6w2, v8r7w1, v9r0w9, v9r1w8, v9r2w7, v9r3w6, v9r4w5,
      v9r5w4, v9r6w3, v9r7w2, vAr0wA, vAr1w9, vAr2w8, vAr3w7,
      vAr4w6, vAr5w5, vAr6w4, vAr7w3, vBr0wB, vBr1wA, vBr2w9,
      vBr3w8, vBr4w7, vBr5w6, vBr6w5, vBr7w4, vCr0wC, vCr1wB,
      vCr2wA, vCr3w9, vCr4w8, vCr5w7, vCr6w6, vCr7w5, vDr0wD,
      vDr1wC, vDr2wB, vDr3wA, vDr4w9, vDr5w8, vDr6w7, vDr7w6,
      vEr0wE, vEr1wD, vEr2wC, vEr3wB, vEr4wA, vEr5w9, vEr6w8,
      vEr7w7, vFr0wF, vFr1wE, vFr2wD, vFr3wC, vFr4wB, vFr5wA,
      vFr6w9, vFr7w8, vGr0wG, vGr1wF, vGr2wE, vGr3wD, vGr4wC,
      vGr5wB, vGr6wA, vGr7w9 );
  end

endmodule
