/****************************************************************
 ---------------------------------------------------------------
     Copyright 1999 Sun Microsystems, Inc., 901 San Antonio
     Road, Palo Alto, CA 94303, U.S.A.  All Rights Reserved.
     The contents of this file are subject to the current
     version of the Sun Community Source License, picoJava-II
     Core ("the License").  You may not use this file except
     in compliance with the License.  You may obtain a copy
     of the License by searching for "Sun Community Source
     License" on the World Wide Web at http://www.sun.com.
     See the License for the rights, obligations, and
     limitations governing use of the contents of this file.

     Sun, Sun Microsystems, the Sun logo, and all Sun-based
     trademarks and logos, Java, picoJava, and all Java-based
     trademarks and logos are trademarks or registered trademarks 
     of Sun Microsystems, Inc. in the United States and other
     countries.
 ----------------------------------------------------------------
******************************************************************/



module mj_s_ff_s_d(out,in, clk);
output out;
input clk;
input in;

reg out;

/* synopsys translate_off */
initial out = 0;
/* synopsys translate_on */

always @(posedge clk)
            out <= #1 in;

endmodule

module mj_s_ff_se_d(out,in, lenable, clk);
output out;
input clk;
input lenable;
input in;
reg out;
always @(posedge clk)
        if (lenable)
            out <= #1 in;
        else
            out <= #1 out;
endmodule

module mj_s_ff_snr_d(out,in, reset_l, clk);
output out;
input clk;
input reset_l;
input in;

reg out;

always @(posedge clk)
        if (~reset_l)
            out <= #1 1'b0;
        else
            out <= #1 in;

endmodule

module mj_s_ff_snre_d(out,in, lenable,reset_l, clk);
output out;
input clk;
input lenable;
input reset_l;
input in;

reg out;
always @(posedge clk)
        if (~reset_l) 
	out <= #1 1'b0;
	else
    	if (lenable)
            out <= #1 in;
        else
            out <= #1 out;

endmodule

/**** Multi Width flops ******/

module mj_s_ff_s_d_2 (out, din, clk);
    output  [1:0]  out;
    input   [1:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]), .clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]), .clk(clk));

endmodule 


module mj_s_ff_se_d_3 (out,din, lenable, clk);
output [2:0] out;
input [2:0] din;
input lenable;
input clk;

mj_s_ff_se_d    mj_s_ff_se_d_0(.out(out[0]),.in(din[0]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_1(.out(out[1]),.in(din[1]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_2(.out(out[2]),.in(din[2]),.lenable(lenable), .clk(clk));

endmodule

module mj_s_ff_se_d_4 (out,din, lenable, clk);
output [3:0] out;
input [3:0] din;
input lenable;
input clk;

mj_s_ff_se_d    mj_s_ff_se_d_0(.out(out[0]),.in(din[0]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_1(.out(out[1]),.in(din[1]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_2(.out(out[2]),.in(din[2]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_3(.out(out[3]),.in(din[3]),.lenable(lenable), .clk(clk));

endmodule

module mj_s_ff_se_d_8 (out,din, lenable, clk);
output [7:0] out;
input [7:0] din;
input lenable;
input clk;

mj_s_ff_se_d    mj_s_ff_se_d_0(.out(out[0]),.in(din[0]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_1(.out(out[1]),.in(din[1]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_2(.out(out[2]),.in(din[2]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_3(.out(out[3]),.in(din[3]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_4(.out(out[4]),.in(din[4]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_5(.out(out[5]),.in(din[5]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_6(.out(out[6]),.in(din[6]),.lenable(lenable), .clk(clk));
mj_s_ff_se_d    mj_s_ff_se_d_7(.out(out[7]),.in(din[7]),.lenable(lenable), .clk(clk));

endmodule

module mj_s_ff_s_d_3 (out, din,clk);
    output  [2:0]  out;
    input   [2:0]  din;
    input           clk; 

mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));

endmodule 


module mj_s_ff_s_d_4 (out, din, clk);
    output  [3:0]  out;
    input   [3:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));

endmodule 


module mj_s_ff_s_d_5 (out, din,clk);
    output  [4:0]  out;
    input   [4:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));

endmodule 


module mj_s_ff_s_d_6 (out, din,clk);
    output  [5:0]  out;
    input   [5:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));

endmodule 


module mj_s_ff_s_d_7 (out, din,clk);
    output  [6:0]  out;
    input   [6:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));

endmodule 


module mj_s_ff_s_d_8 (out, din,clk);
    output  [7:0]  out;
    input   [7:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));   
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));

endmodule 


module mj_s_ff_s_d_9 (out, din,clk);
    output  [8:0]  out;
    input   [8:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));

endmodule 


module mj_s_ff_s_d_10 (out, din,clk);
    output  [9:0]  out;
    input   [9:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));


endmodule 


module mj_s_ff_s_d_11 (out, din,clk);
    output  [10:0]  out;
    input   [10:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));

        

endmodule 


module mj_s_ff_s_d_12 (out, din,clk);
    output  [11:0]  out;
    input   [11:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
 
endmodule 

module mj_s_ff_s_d_13 (out, din,clk);
    output  [12:0]  out;
    input   [12:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
    
endmodule 

module mj_s_ff_s_d_14 (out, din,clk);
    output  [13:0]  out;
    input   [13:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));

endmodule 

module mj_s_ff_s_d_15 (out, din,clk);
    output  [14:0]  out;
    input   [14:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
   
endmodule 

module mj_s_ff_s_d_16 (out, din,clk);
    output  [15:0]  out;
    input   [15:0]  din;
    input           clk;

mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));

endmodule 

module mj_s_ff_s_d_17 (out, din,clk);
    output  [16:0]  out;
    input   [16:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));

    
endmodule 


module mj_s_ff_s_d_18 (out, din,clk);
    output  [17:0]  out;
    input   [17:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));

endmodule 


module mj_s_ff_s_d_19 (out, din,clk);
    output  [18:0]  out;
    input   [18:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));   
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));


endmodule 


module mj_s_ff_s_d_20 (out, din,clk);
    output  [19:0]  out;
    input   [19:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));


endmodule 


module mj_s_ff_s_d_21 (out, din,clk);
    output  [20:0]  out;
    input   [20:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));

endmodule 


module mj_s_ff_s_d_22 (out, din,clk);
    output  [21:0]  out;
    input   [21:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));


    
endmodule 


module mj_s_ff_s_d_23 (out, din,clk);
    output  [22:0]  out;
    input   [22:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));

  
endmodule 


module mj_s_ff_s_d_24 (out, din,clk);
    output  [23:0]  out;
    input   [23:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));

   
endmodule 


module mj_s_ff_s_d_25 (out, din,clk);
    output  [24:0]  out;
    input   [24:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));

  
endmodule 


module mj_s_ff_s_d_26 (out, din,clk);
    output  [25:0]  out;
    input   [25:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));


   endmodule 


module mj_s_ff_s_d_27 (out, din,clk);
    output  [26:0]  out;
    input   [26:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.clk(clk));

endmodule 

module mj_s_ff_s_d_28 (out, din,clk);
    output  [27:0]  out;
    input   [27:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_27(.out(out[27]),.in(din[27]),.clk(clk));

  
endmodule 


module mj_s_ff_s_d_29 (out, din,clk);
    output  [28:0]  out;
    input   [28:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_27(.out(out[27]),.in(din[27]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_28(.out(out[28]),.in(din[28]),.clk(clk));

endmodule 


module mj_s_ff_s_d_30 (out, din,clk);
    output  [29:0]  out;
    input   [29:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_27(.out(out[27]),.in(din[27]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_28(.out(out[28]),.in(din[28]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_29(.out(out[29]),.in(din[29]),.clk(clk));


endmodule 


module mj_s_ff_s_d_31 (out, din,clk);
    output  [30:0]  out;
    input   [30:0]  din;
    input           clk;
mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));    
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_27(.out(out[27]),.in(din[27]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_28(.out(out[28]),.in(din[28]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_29(.out(out[29]),.in(din[29]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_30(.out(out[30]),.in(din[30]),.clk(clk));

endmodule 

module mj_s_ff_se_d_32 (out,din, lenable,clk);
output [31:0] out;
input clk;
input lenable;
input [31:0] din;

mj_s_ff_se_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_27(.out(out[27]),.in(din[27]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_28(.out(out[28]),.in(din[28]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_29(.out(out[29]),.in(din[29]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_30(.out(out[30]),.in(din[30]),.lenable(lenable),.clk(clk));
mj_s_ff_se_d    mj_s_ff_s_d_31(.out(out[31]),.in(din[31]),.lenable(lenable),.clk(clk));

endmodule

module mj_s_ff_s_d_32 (out, din,clk);
    output  [31:0]  out;
    input   [31:0]  din;
    input           clk; 

mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(din[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(din[1]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(din[2]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(din[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(din[4]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(din[5]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(din[6]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(din[7]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(din[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(din[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(din[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(din[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(din[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(din[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(din[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(din[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(din[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(din[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(din[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(din[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(din[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(din[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(din[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(din[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(din[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(din[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(din[26]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_27(.out(out[27]),.in(din[27]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_28(.out(out[28]),.in(din[28]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_29(.out(out[29]),.in(din[29]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_30(.out(out[30]),.in(din[30]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_31(.out(out[31]),.in(din[31]),.clk(clk));

endmodule 

module mj_s_ff_snr_d_2 (out, din, reset_l,clk);
    output  [1:0]  out;
    input   [1:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_3 (out, din, reset_l,clk);
    output  [2:0]  out;
    input   [2:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_4 (out, din, reset_l,clk);
    output  [3:0]  out;
    input   [3:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_5 (out, din, reset_l,clk);
    output  [4:0]  out;
    input   [4:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_6 (out, din, reset_l,clk);
    output  [5:0]  out;
    input   [5:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_7 (out, din, reset_l,clk);
    output  [6:0]  out;
    input   [6:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_8 (out, din, reset_l,clk);
    output  [7:0]  out;
    input   [7:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_9 (out, din, reset_l,clk);
    output  [8:0]  out;
    input   [8:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_10 (out, din, reset_l,clk);
    output  [9:0]  out;
    input   [9:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_11 (out, din, reset_l,clk);
    output  [10:0]  out;
    input   [10:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_12 (out, din, reset_l,clk);
    output  [11:0]  out;
    input   [11:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_13 (out, din, reset_l,clk);
    output  [12:0]  out;
    input   [12:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_14 (out, din, reset_l,clk);
    output  [13:0]  out;
    input   [13:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_15 (out, din, reset_l,clk);
    output  [14:0]  out;
    input   [14:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_16 (out, din, reset_l,clk);
    output  [15:0]  out;
    input   [15:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_17 (out, din, reset_l,clk);
    output  [16:0]  out;
    input   [16:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_18 (out, din, reset_l,clk);
    output  [17:0]  out;
    input   [17:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_19 (out, din, reset_l,clk);
    output  [18:0]  out;
    input   [18:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_20 (out, din, reset_l,clk);
    output  [19:0]  out;
    input   [19:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_21 (out, din, reset_l,clk);
    output  [20:0]  out;
    input   [20:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_22 (out, din, reset_l,clk);
    output  [21:0]  out;
    input   [21:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_23 (out, din, reset_l,clk);
    output  [22:0]  out;
    input   [22:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_24 (out, din, reset_l,clk);
    output  [23:0]  out;
    input   [23:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_25 (out, din, reset_l,clk);
    output  [24:0]  out;
    input   [24:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_26 (out, din, reset_l,clk);
    output  [25:0]  out;
    input   [25:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_27 (out, din, reset_l,clk);
    output  [26:0]  out;
    input   [26:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_28 (out, din, reset_l,clk);
    output  [27:0]  out;
    input   [27:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_27(.out(out[27]), .in(din[27]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_29 (out, din, reset_l,clk);
    output  [28:0]  out;
    input   [28:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_27(.out(out[27]), .in(din[27]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_28(.out(out[28]), .in(din[28]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_30 (out, din, reset_l,clk);
    output  [29:0]  out;
    input   [29:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_27(.out(out[27]), .in(din[27]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_28(.out(out[28]), .in(din[28]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_29(.out(out[29]), .in(din[29]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_31 (out, din, reset_l,clk);
    output  [30:0]  out;
    input   [30:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_27(.out(out[27]), .in(din[27]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_28(.out(out[28]), .in(din[28]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_29(.out(out[29]), .in(din[29]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_30(.out(out[30]), .in(din[30]), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_32 (out, din, reset_l,clk);
    output  [31:0]  out;
    input   [31:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_27(.out(out[27]), .in(din[27]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_28(.out(out[28]), .in(din[28]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_29(.out(out[29]), .in(din[29]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_30(.out(out[30]), .in(din[30]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_31(.out(out[31]), .in(din[31]), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_6 (out, din, lenable, reset_l,clk);
    output  [5:0]  out;
    input   [5:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;
 
    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
 
endmodule

module mj_s_ff_snre_d_7 (out, din, lenable, reset_l,clk);
    output  [6:0]  out;
    input   [6:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;
 
    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
 
endmodule

module mj_s_ff_snre_d_8 (out, din, lenable, reset_l,clk);
    output  [7:0]  out;
    input   [7:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_12 (out, din, lenable, reset_l,clk);
    output  [11:0]  out;
    input   [11:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_16 (out, din, lenable, reset_l,clk);
    output  [15:0]  out;
    input   [15:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_23 (out, din, lenable, reset_l,clk);
    output  [22:0]  out;
    input   [22:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snre_d_30 (out, din, lenable, reset_l,clk);
    output  [29:0]  out;
    input   [29:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_23(.out(out[23]), .in(din[23]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_24(.out(out[24]), .in(din[24]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_25(.out(out[25]), .in(din[25]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_26(.out(out[26]), .in(din[26]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_27(.out(out[27]), .in(din[27]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_28(.out(out[28]), .in(din[28]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_29(.out(out[29]), .in(din[29]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_32 (out, din, lenable, reset_l,clk);
    output  [31:0]  out;
    input   [31:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_23(.out(out[23]), .in(din[23]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_24(.out(out[24]), .in(din[24]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_25(.out(out[25]), .in(din[25]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_26(.out(out[26]), .in(din[26]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_27(.out(out[27]), .in(din[27]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_28(.out(out[28]), .in(din[28]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_29(.out(out[29]), .in(din[29]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_30(.out(out[30]), .in(din[30]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_31(.out(out[31]), .in(din[31]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snr_d_64 (out, din, reset_l,clk);
    output  [63:0]  out;
    input   [63:0]  din;
    input           clk;
    input           reset_l;

    mj_s_ff_snr_d    mj_s_ff_snr_d_0(.out(out[0]), .in(din[0]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_1(.out(out[1]), .in(din[1]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_2(.out(out[2]), .in(din[2]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_3(.out(out[3]), .in(din[3]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_4(.out(out[4]), .in(din[4]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_5(.out(out[5]), .in(din[5]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_6(.out(out[6]), .in(din[6]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_7(.out(out[7]), .in(din[7]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_8(.out(out[8]), .in(din[8]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_9(.out(out[9]), .in(din[9]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_10(.out(out[10]), .in(din[10]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_11(.out(out[11]), .in(din[11]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_12(.out(out[12]), .in(din[12]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_13(.out(out[13]), .in(din[13]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_14(.out(out[14]), .in(din[14]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_15(.out(out[15]), .in(din[15]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_16(.out(out[16]), .in(din[16]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_17(.out(out[17]), .in(din[17]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_18(.out(out[18]), .in(din[18]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_19(.out(out[19]), .in(din[19]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_20(.out(out[20]), .in(din[20]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_21(.out(out[21]), .in(din[21]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_22(.out(out[22]), .in(din[22]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_23(.out(out[23]), .in(din[23]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_24(.out(out[24]), .in(din[24]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_25(.out(out[25]), .in(din[25]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_26(.out(out[26]), .in(din[26]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_27(.out(out[27]), .in(din[27]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_28(.out(out[28]), .in(din[28]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_29(.out(out[29]), .in(din[29]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_30(.out(out[30]), .in(din[30]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_31(.out(out[31]), .in(din[31]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_32(.out(out[32]), .in(din[32]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_33(.out(out[33]), .in(din[33]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_34(.out(out[34]), .in(din[34]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_35(.out(out[35]), .in(din[35]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_36(.out(out[36]), .in(din[36]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_37(.out(out[37]), .in(din[37]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_38(.out(out[38]), .in(din[38]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_39(.out(out[39]), .in(din[39]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_40(.out(out[40]), .in(din[40]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_41(.out(out[41]), .in(din[41]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_42(.out(out[42]), .in(din[42]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_43(.out(out[43]), .in(din[43]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_44(.out(out[44]), .in(din[44]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_45(.out(out[45]), .in(din[45]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_46(.out(out[46]), .in(din[46]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_47(.out(out[47]), .in(din[47]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_48(.out(out[48]), .in(din[48]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_49(.out(out[49]), .in(din[49]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_50(.out(out[50]), .in(din[50]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_51(.out(out[51]), .in(din[51]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_52(.out(out[52]), .in(din[52]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_53(.out(out[53]), .in(din[53]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_54(.out(out[54]), .in(din[54]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_55(.out(out[55]), .in(din[55]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_56(.out(out[56]), .in(din[56]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_57(.out(out[57]), .in(din[57]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_58(.out(out[58]), .in(din[58]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_59(.out(out[59]), .in(din[59]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_60(.out(out[60]), .in(din[60]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_61(.out(out[61]), .in(din[61]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_62(.out(out[62]), .in(din[62]), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snr_d    mj_s_ff_snr_d_63(.out(out[63]), .in(din[63]), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_s_d_64 (out, in, clk);
output  [63:0]  out;
input           clk;
input   [63:0]  in;

wire    [63:0]  out;

mj_s_ff_s_d    mj_s_ff_s_d_0(.out(out[0]),.in(in[0]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_1(.out(out[1]),.in(in[1]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_2(.out(out[2]),.in(in[2]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_3(.out(out[3]),.in(in[3]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_4(.out(out[4]),.in(in[4]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_5(.out(out[5]),.in(in[5]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_6(.out(out[6]),.in(in[6]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_7(.out(out[7]),.in(in[7]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_8(.out(out[8]),.in(in[8]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_9(.out(out[9]),.in(in[9]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_10(.out(out[10]),.in(in[10]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_11(.out(out[11]),.in(in[11]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_12(.out(out[12]),.in(in[12]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_13(.out(out[13]),.in(in[13]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_14(.out(out[14]),.in(in[14]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_15(.out(out[15]),.in(in[15]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_16(.out(out[16]),.in(in[16]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_17(.out(out[17]),.in(in[17]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_18(.out(out[18]),.in(in[18]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_19(.out(out[19]),.in(in[19]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_20(.out(out[20]),.in(in[20]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_21(.out(out[21]),.in(in[21]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_22(.out(out[22]),.in(in[22]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_23(.out(out[23]),.in(in[23]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_24(.out(out[24]),.in(in[24]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_25(.out(out[25]),.in(in[25]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_26(.out(out[26]),.in(in[26]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_27(.out(out[27]),.in(in[27]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_28(.out(out[28]),.in(in[28]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_29(.out(out[29]),.in(in[29]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_30(.out(out[30]),.in(in[30]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_31(.out(out[31]),.in(in[31]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_32(.out(out[32]),.in(in[32]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_33(.out(out[33]),.in(in[33]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_34(.out(out[34]),.in(in[34]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_35(.out(out[35]),.in(in[35]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_36(.out(out[36]),.in(in[36]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_37(.out(out[37]),.in(in[37]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_38(.out(out[38]),.in(in[38]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_39(.out(out[39]),.in(in[39]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_40(.out(out[40]),.in(in[40]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_41(.out(out[41]),.in(in[41]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_42(.out(out[42]),.in(in[42]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_43(.out(out[43]),.in(in[43]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_44(.out(out[44]),.in(in[44]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_45(.out(out[45]),.in(in[45]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_46(.out(out[46]),.in(in[46]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_47(.out(out[47]),.in(in[47]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_48(.out(out[48]),.in(in[48]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_49(.out(out[49]),.in(in[49]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_50(.out(out[50]),.in(in[50]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_51(.out(out[51]),.in(in[51]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_52(.out(out[52]),.in(in[52]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_53(.out(out[53]),.in(in[53]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_54(.out(out[54]),.in(in[54]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_55(.out(out[55]),.in(in[55]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_56(.out(out[56]),.in(in[56]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_57(.out(out[57]),.in(in[57]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_58(.out(out[58]),.in(in[58]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_59(.out(out[59]),.in(in[59]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_60(.out(out[60]),.in(in[60]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_61(.out(out[61]),.in(in[61]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_62(.out(out[62]),.in(in[62]),.clk(clk));
mj_s_ff_s_d    mj_s_ff_s_d_63(.out(out[63]),.in(in[63]),.clk(clk));
endmodule




module ff_s (out, din, clk) ;
    output    out;
    input     din;
    input     clk;
 
mj_s_ff_s_d  mj_s_ff_s_d_0 (	.out(out),
				.in(din),
				.clk(clk)
				);
endmodule


module ff_sre(out, din, enable, reset_l, clk) ;
    output   out;
    input    din;
    input    clk;
    input    reset_l;
    input    enable;
 
mj_s_ff_snre_d  mj_s_ff_snre_d_0 (      .out(out),
                                        .in(din), 
                                        .lenable(enable),
                                        .reset_l(reset_l),
                                        .clk(clk)
                                        );
endmodule


module ff_se (out, din, enable, clk) ;
    output    out;
    input     din;
    input     clk;
    input     enable;
 
mj_s_ff_se_d  mj_s_ff_se_d_0 (  .out(out),
                                .in(din),
                                .lenable(enable),
                                .clk(clk)
                                );

endmodule


module ff_sr(out, din, reset_l, clk) ;
    output   out;
    input    din;
    input    clk;
    input    reset_l;
 
mj_s_ff_snr_d  mj_s_ff_snr_d_0 (        .out(out),
                                        .in(din),
                                        .reset_l(reset_l),
                                        .clk(clk)
                                        );
endmodule



module ff_s_2 (out, din, clk) ;
    output  [1:0]  out;
    input   [1:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);

endmodule 


module ff_s_3 (out, din, clk) ;
    output  [2:0]  out;
    input   [2:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);

endmodule 


module ff_s_4 (out, din, clk) ;
    output  [3:0]  out;
    input   [3:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);

endmodule 


module ff_s_5 (out, din, clk) ;
    output  [4:0]  out;
    input   [4:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);

endmodule 


module ff_s_6 (out, din, clk) ;
    output  [5:0]  out;
    input   [5:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);

endmodule 


module ff_s_7 (out, din, clk) ;
    output  [6:0]  out;
    input   [6:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);

endmodule 


module ff_s_8 (out, din, clk) ;
    output  [7:0]  out;
    input   [7:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);

endmodule 


module ff_s_9 (out, din, clk) ;
    output  [8:0]  out;
    input   [8:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);

endmodule 


module ff_s_10 (out, din, clk) ;
    output  [9:0]  out;
    input   [9:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);

endmodule 


module ff_s_11 (out, din, clk) ;
    output  [10:0]  out;
    input   [10:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);

endmodule 


module ff_s_12 (out, din, clk) ;
    output  [11:0]  out;
    input   [11:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);

endmodule 


module ff_s_13 (out, din, clk) ;
    output  [12:0]  out;
    input   [12:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);

endmodule 


module ff_s_14 (out, din, clk) ;
    output  [13:0]  out;
    input   [13:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);

endmodule 


module ff_s_15 (out, din, clk) ;
    output  [14:0]  out;
    input   [14:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);

endmodule 


module ff_s_16 (out, din, clk) ;
    output  [15:0]  out;
    input   [15:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);

endmodule 


module ff_s_17 (out, din, clk) ;
    output  [16:0]  out;
    input   [16:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);

endmodule 


module ff_s_18 (out, din, clk) ;
    output  [17:0]  out;
    input   [17:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);

endmodule 


module ff_s_19 (out, din, clk) ;
    output  [18:0]  out;
    input   [18:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);

endmodule 


module ff_s_20 (out, din, clk) ;
    output  [19:0]  out;
    input   [19:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);

endmodule 


module ff_s_21 (out, din, clk) ;
    output  [20:0]  out;
    input   [20:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);

endmodule 


module ff_s_22 (out, din, clk) ;
    output  [21:0]  out;
    input   [21:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);

endmodule 


module ff_s_23 (out, din, clk) ;
    output  [22:0]  out;
    input   [22:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);

endmodule 


module ff_s_24 (out, din, clk) ;
    output  [23:0]  out;
    input   [23:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);

endmodule 


module ff_s_25 (out, din, clk) ;
    output  [24:0]  out;
    input   [24:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);

endmodule 


module ff_s_26 (out, din, clk) ;
    output  [25:0]  out;
    input   [25:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);

endmodule 


module ff_s_27 (out, din, clk) ;
    output  [26:0]  out;
    input   [26:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);

endmodule 


module ff_s_28 (out, din, clk) ;
    output  [27:0]  out;
    input   [27:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);
    ff_s    ff_s_27(out[27], din[27], clk);

endmodule 


module ff_s_29 (out, din, clk) ;
    output  [28:0]  out;
    input   [28:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);
    ff_s    ff_s_27(out[27], din[27], clk);
    ff_s    ff_s_28(out[28], din[28], clk);

endmodule 


module ff_s_30 (out, din, clk) ;
    output  [29:0]  out;
    input   [29:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);
    ff_s    ff_s_27(out[27], din[27], clk);
    ff_s    ff_s_28(out[28], din[28], clk);
    ff_s    ff_s_29(out[29], din[29], clk);

endmodule 


module ff_s_31 (out, din, clk) ;
    output  [30:0]  out;
    input   [30:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);
    ff_s    ff_s_27(out[27], din[27], clk);
    ff_s    ff_s_28(out[28], din[28], clk);
    ff_s    ff_s_29(out[29], din[29], clk);
    ff_s    ff_s_30(out[30], din[30], clk);

endmodule 


module ff_s_32 (out, din, clk) ;
    output  [31:0]  out;
    input   [31:0]  din;
    input           clk;

    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);
    ff_s    ff_s_27(out[27], din[27], clk);
    ff_s    ff_s_28(out[28], din[28], clk);
    ff_s    ff_s_29(out[29], din[29], clk);
    ff_s    ff_s_30(out[30], din[30], clk);
    ff_s    ff_s_31(out[31], din[31], clk);

endmodule 


module ff_se_2 (out, din, enable, clk) ;
    output  [1:0]  out;
    input   [1:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);

endmodule 


module ff_se_3 (out, din, enable, clk) ;
    output  [2:0]  out;
    input   [2:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);

endmodule 


module ff_se_4 (out, din, enable, clk) ;
    output  [3:0]  out;
    input   [3:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);

endmodule 


module ff_se_5 (out, din, enable, clk) ;
    output  [4:0]  out;
    input   [4:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);

endmodule 


module ff_se_6 (out, din, enable, clk) ;
    output  [5:0]  out;
    input   [5:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);

endmodule 


module ff_se_7 (out, din, enable, clk) ;
    output  [6:0]  out;
    input   [6:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);

endmodule 


module ff_se_8 (out, din, enable, clk) ;
    output  [7:0]  out;
    input   [7:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);

endmodule 


module ff_se_9 (out, din, enable, clk) ;
    output  [8:0]  out;
    input   [8:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);

endmodule 


module ff_se_10 (out, din, enable, clk) ;
    output  [9:0]  out;
    input   [9:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);

endmodule 


module ff_se_11 (out, din, enable, clk) ;
    output  [10:0]  out;
    input   [10:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);

endmodule 


module ff_se_12 (out, din, enable, clk) ;
    output  [11:0]  out;
    input   [11:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);

endmodule 


module ff_se_13 (out, din, enable, clk) ;
    output  [12:0]  out;
    input   [12:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);

endmodule 


module ff_se_14 (out, din, enable, clk) ;
    output  [13:0]  out;
    input   [13:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);

endmodule 


module ff_se_15 (out, din, enable, clk) ;
    output  [14:0]  out;
    input   [14:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);

endmodule 


module ff_se_16 (out, din, enable, clk) ;
    output  [15:0]  out;
    input   [15:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);

endmodule 


module ff_se_17 (out, din, enable, clk) ;
    output  [16:0]  out;
    input   [16:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);

endmodule 


module ff_se_18 (out, din, enable, clk) ;
    output  [17:0]  out;
    input   [17:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);

endmodule 


module ff_se_19 (out, din, enable, clk) ;
    output  [18:0]  out;
    input   [18:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);

endmodule 


module ff_se_20 (out, din, enable, clk) ;
    output  [19:0]  out;
    input   [19:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);

endmodule 


module ff_se_21 (out, din, enable, clk) ;
    output  [20:0]  out;
    input   [20:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);

endmodule 


module ff_se_22 (out, din, enable, clk) ;
    output  [21:0]  out;
    input   [21:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);

endmodule 


module ff_se_23 (out, din, enable, clk) ;
    output  [22:0]  out;
    input   [22:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);

endmodule 


module ff_se_24 (out, din, enable, clk) ;
    output  [23:0]  out;
    input   [23:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);

endmodule 


module ff_se_25 (out, din, enable, clk) ;
    output  [24:0]  out;
    input   [24:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);

endmodule 


module ff_se_26 (out, din, enable, clk) ;
    output  [25:0]  out;
    input   [25:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);

endmodule 


module ff_se_27 (out, din, enable, clk) ;
    output  [26:0]  out;
    input   [26:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);
    ff_se    ff_se_26(out[26], din[26], enable, clk);

endmodule 


module ff_se_28 (out, din, enable, clk) ;
    output  [27:0]  out;
    input   [27:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);
    ff_se    ff_se_26(out[26], din[26], enable, clk);
    ff_se    ff_se_27(out[27], din[27], enable, clk);

endmodule 


module ff_se_29 (out, din, enable, clk) ;
    output  [28:0]  out;
    input   [28:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);
    ff_se    ff_se_26(out[26], din[26], enable, clk);
    ff_se    ff_se_27(out[27], din[27], enable, clk);
    ff_se    ff_se_28(out[28], din[28], enable, clk);

endmodule 


module ff_se_30 (out, din, enable, clk) ;
    output  [29:0]  out;
    input   [29:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);
    ff_se    ff_se_26(out[26], din[26], enable, clk);
    ff_se    ff_se_27(out[27], din[27], enable, clk);
    ff_se    ff_se_28(out[28], din[28], enable, clk);
    ff_se    ff_se_29(out[29], din[29], enable, clk);

endmodule 


module ff_se_31 (out, din, enable, clk) ;
    output  [30:0]  out;
    input   [30:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);
    ff_se    ff_se_26(out[26], din[26], enable, clk);
    ff_se    ff_se_27(out[27], din[27], enable, clk);
    ff_se    ff_se_28(out[28], din[28], enable, clk);
    ff_se    ff_se_29(out[29], din[29], enable, clk);
    ff_se    ff_se_30(out[30], din[30], enable, clk);

endmodule 


module ff_se_32 (out, din, enable, clk) ;
    output  [31:0]  out;
    input   [31:0]  din;
    input           clk;
    input           enable;

    ff_se    ff_se_0(out[0], din[0], enable, clk);
    ff_se    ff_se_1(out[1], din[1], enable, clk);
    ff_se    ff_se_2(out[2], din[2], enable, clk);
    ff_se    ff_se_3(out[3], din[3], enable, clk);
    ff_se    ff_se_4(out[4], din[4], enable, clk);
    ff_se    ff_se_5(out[5], din[5], enable, clk);
    ff_se    ff_se_6(out[6], din[6], enable, clk);
    ff_se    ff_se_7(out[7], din[7], enable, clk);
    ff_se    ff_se_8(out[8], din[8], enable, clk);
    ff_se    ff_se_9(out[9], din[9], enable, clk);
    ff_se    ff_se_10(out[10], din[10], enable, clk);
    ff_se    ff_se_11(out[11], din[11], enable, clk);
    ff_se    ff_se_12(out[12], din[12], enable, clk);
    ff_se    ff_se_13(out[13], din[13], enable, clk);
    ff_se    ff_se_14(out[14], din[14], enable, clk);
    ff_se    ff_se_15(out[15], din[15], enable, clk);
    ff_se    ff_se_16(out[16], din[16], enable, clk);
    ff_se    ff_se_17(out[17], din[17], enable, clk);
    ff_se    ff_se_18(out[18], din[18], enable, clk);
    ff_se    ff_se_19(out[19], din[19], enable, clk);
    ff_se    ff_se_20(out[20], din[20], enable, clk);
    ff_se    ff_se_21(out[21], din[21], enable, clk);
    ff_se    ff_se_22(out[22], din[22], enable, clk);
    ff_se    ff_se_23(out[23], din[23], enable, clk);
    ff_se    ff_se_24(out[24], din[24], enable, clk);
    ff_se    ff_se_25(out[25], din[25], enable, clk);
    ff_se    ff_se_26(out[26], din[26], enable, clk);
    ff_se    ff_se_27(out[27], din[27], enable, clk);
    ff_se    ff_se_28(out[28], din[28], enable, clk);
    ff_se    ff_se_29(out[29], din[29], enable, clk);
    ff_se    ff_se_30(out[30], din[30], enable, clk);
    ff_se    ff_se_31(out[31], din[31], enable, clk);

endmodule 


module ff_sr_2 (out, din, reset_l, clk) ;
    output  [1:0]  out;
    input   [1:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);

endmodule 


module ff_sr_3 (out, din, reset_l, clk) ;
    output  [2:0]  out;
    input   [2:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);

endmodule 


module ff_sr_4 (out, din, reset_l, clk) ;
    output  [3:0]  out;
    input   [3:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);

endmodule 


module ff_sr_5 (out, din, reset_l, clk) ;
    output  [4:0]  out;
    input   [4:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);

endmodule 


module ff_sr_6 (out, din, reset_l, clk) ;
    output  [5:0]  out;
    input   [5:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);

endmodule 


module ff_sr_7 (out, din, reset_l, clk) ;
    output  [6:0]  out;
    input   [6:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);

endmodule 


module ff_sr_8 (out, din, reset_l, clk) ;
    output  [7:0]  out;
    input   [7:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);

endmodule 


module ff_sr_9 (out, din, reset_l, clk) ;
    output  [8:0]  out;
    input   [8:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);

endmodule 


module ff_sr_10 (out, din, reset_l, clk) ;
    output  [9:0]  out;
    input   [9:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);

endmodule 


module ff_sr_11 (out, din, reset_l, clk) ;
    output  [10:0]  out;
    input   [10:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);

endmodule 


module ff_sr_12 (out, din, reset_l, clk) ;
    output  [11:0]  out;
    input   [11:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);

endmodule 


module ff_sr_13 (out, din, reset_l, clk) ;
    output  [12:0]  out;
    input   [12:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);

endmodule 


module ff_sr_14 (out, din, reset_l, clk) ;
    output  [13:0]  out;
    input   [13:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);

endmodule 


module ff_sr_15 (out, din, reset_l, clk) ;
    output  [14:0]  out;
    input   [14:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);

endmodule 


module ff_sr_16 (out, din, reset_l, clk) ;
    output  [15:0]  out;
    input   [15:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);

endmodule 


module ff_sr_17 (out, din, reset_l, clk) ;
    output  [16:0]  out;
    input   [16:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);

endmodule 


module ff_sr_18 (out, din, reset_l, clk) ;
    output  [17:0]  out;
    input   [17:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);

endmodule 


module ff_sr_19 (out, din, reset_l, clk) ;
    output  [18:0]  out;
    input   [18:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);

endmodule 


module ff_sr_20 (out, din, reset_l, clk) ;
    output  [19:0]  out;
    input   [19:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);

endmodule 


module ff_sr_21 (out, din, reset_l, clk) ;
    output  [20:0]  out;
    input   [20:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);

endmodule 


module ff_sr_22 (out, din, reset_l, clk) ;
    output  [21:0]  out;
    input   [21:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);

endmodule 


module ff_sr_23 (out, din, reset_l, clk) ;
    output  [22:0]  out;
    input   [22:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);

endmodule 


module ff_sr_24 (out, din, reset_l, clk) ;
    output  [23:0]  out;
    input   [23:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);

endmodule 


module ff_sr_25 (out, din, reset_l, clk) ;
    output  [24:0]  out;
    input   [24:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);

endmodule 


module ff_sr_26 (out, din, reset_l, clk) ;
    output  [25:0]  out;
    input   [25:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);

endmodule 


module ff_sr_27 (out, din, reset_l, clk) ;
    output  [26:0]  out;
    input   [26:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);
    ff_sr    ff_sr_26(out[26], din[26], reset_l, clk);

endmodule 


module ff_sr_28 (out, din, reset_l, clk) ;
    output  [27:0]  out;
    input   [27:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);
    ff_sr    ff_sr_26(out[26], din[26], reset_l, clk);
    ff_sr    ff_sr_27(out[27], din[27], reset_l, clk);

endmodule 


module ff_sr_29 (out, din, reset_l, clk) ;
    output  [28:0]  out;
    input   [28:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);
    ff_sr    ff_sr_26(out[26], din[26], reset_l, clk);
    ff_sr    ff_sr_27(out[27], din[27], reset_l, clk);
    ff_sr    ff_sr_28(out[28], din[28], reset_l, clk);

endmodule 


module ff_sr_30 (out, din, reset_l, clk) ;
    output  [29:0]  out;
    input   [29:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);
    ff_sr    ff_sr_26(out[26], din[26], reset_l, clk);
    ff_sr    ff_sr_27(out[27], din[27], reset_l, clk);
    ff_sr    ff_sr_28(out[28], din[28], reset_l, clk);
    ff_sr    ff_sr_29(out[29], din[29], reset_l, clk);

endmodule 


module ff_sr_31 (out, din, reset_l, clk) ;
    output  [30:0]  out;
    input   [30:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);
    ff_sr    ff_sr_26(out[26], din[26], reset_l, clk);
    ff_sr    ff_sr_27(out[27], din[27], reset_l, clk);
    ff_sr    ff_sr_28(out[28], din[28], reset_l, clk);
    ff_sr    ff_sr_29(out[29], din[29], reset_l, clk);
    ff_sr    ff_sr_30(out[30], din[30], reset_l, clk);

endmodule 


module ff_sr_32 (out, din, reset_l, clk) ;
    output  [31:0]  out;
    input   [31:0]  din;
    input           clk;
    input           reset_l;

    ff_sr    ff_sr_0(out[0], din[0], reset_l, clk);
    ff_sr    ff_sr_1(out[1], din[1], reset_l, clk);
    ff_sr    ff_sr_2(out[2], din[2], reset_l, clk);
    ff_sr    ff_sr_3(out[3], din[3], reset_l, clk);
    ff_sr    ff_sr_4(out[4], din[4], reset_l, clk);
    ff_sr    ff_sr_5(out[5], din[5], reset_l, clk);
    ff_sr    ff_sr_6(out[6], din[6], reset_l, clk);
    ff_sr    ff_sr_7(out[7], din[7], reset_l, clk);
    ff_sr    ff_sr_8(out[8], din[8], reset_l, clk);
    ff_sr    ff_sr_9(out[9], din[9], reset_l, clk);
    ff_sr    ff_sr_10(out[10], din[10], reset_l, clk);
    ff_sr    ff_sr_11(out[11], din[11], reset_l, clk);
    ff_sr    ff_sr_12(out[12], din[12], reset_l, clk);
    ff_sr    ff_sr_13(out[13], din[13], reset_l, clk);
    ff_sr    ff_sr_14(out[14], din[14], reset_l, clk);
    ff_sr    ff_sr_15(out[15], din[15], reset_l, clk);
    ff_sr    ff_sr_16(out[16], din[16], reset_l, clk);
    ff_sr    ff_sr_17(out[17], din[17], reset_l, clk);
    ff_sr    ff_sr_18(out[18], din[18], reset_l, clk);
    ff_sr    ff_sr_19(out[19], din[19], reset_l, clk);
    ff_sr    ff_sr_20(out[20], din[20], reset_l, clk);
    ff_sr    ff_sr_21(out[21], din[21], reset_l, clk);
    ff_sr    ff_sr_22(out[22], din[22], reset_l, clk);
    ff_sr    ff_sr_23(out[23], din[23], reset_l, clk);
    ff_sr    ff_sr_24(out[24], din[24], reset_l, clk);
    ff_sr    ff_sr_25(out[25], din[25], reset_l, clk);
    ff_sr    ff_sr_26(out[26], din[26], reset_l, clk);
    ff_sr    ff_sr_27(out[27], din[27], reset_l, clk);
    ff_sr    ff_sr_28(out[28], din[28], reset_l, clk);
    ff_sr    ff_sr_29(out[29], din[29], reset_l, clk);
    ff_sr    ff_sr_30(out[30], din[30], reset_l, clk);
    ff_sr    ff_sr_31(out[31], din[31], reset_l, clk);

endmodule 


module ff_sre_2 (out, din, enable, reset_l, clk) ;
    output  [1:0]  out;
    input   [1:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);

endmodule 


module ff_sre_3 (out, din, enable, reset_l, clk) ;
    output  [2:0]  out;
    input   [2:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);

endmodule 


module ff_sre_4 (out, din, enable, reset_l, clk) ;
    output  [3:0]  out;
    input   [3:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);

endmodule 


module ff_sre_5 (out, din, enable, reset_l, clk) ;
    output  [4:0]  out;
    input   [4:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);

endmodule 


module ff_sre_6 (out, din, enable, reset_l, clk) ;
    output  [5:0]  out;
    input   [5:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);

endmodule 


module ff_sre_7 (out, din, enable, reset_l, clk) ;
    output  [6:0]  out;
    input   [6:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);

endmodule 


module ff_sre_8 (out, din, enable, reset_l, clk) ;
    output  [7:0]  out;
    input   [7:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);

endmodule 


module ff_sre_9 (out, din, enable, reset_l, clk) ;
    output  [8:0]  out;
    input   [8:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);

endmodule 


module ff_sre_10 (out, din, enable, reset_l, clk) ;
    output  [9:0]  out;
    input   [9:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);

endmodule 


module ff_sre_11 (out, din, enable, reset_l, clk) ;
    output  [10:0]  out;
    input   [10:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);

endmodule 


module ff_sre_12 (out, din, enable, reset_l, clk) ;
    output  [11:0]  out;
    input   [11:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);

endmodule 


module ff_sre_13 (out, din, enable, reset_l, clk) ;
    output  [12:0]  out;
    input   [12:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);

endmodule 


module ff_sre_14 (out, din, enable, reset_l, clk) ;
    output  [13:0]  out;
    input   [13:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);

endmodule 


module ff_sre_15 (out, din, enable, reset_l, clk) ;
    output  [14:0]  out;
    input   [14:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);

endmodule 


module ff_sre_16 (out, din, enable, reset_l, clk) ;
    output  [15:0]  out;
    input   [15:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);

endmodule 


module ff_sre_17 (out, din, enable, reset_l, clk) ;
    output  [16:0]  out;
    input   [16:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);

endmodule 


module ff_sre_18 (out, din, enable, reset_l, clk) ;
    output  [17:0]  out;
    input   [17:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);

endmodule 


module ff_sre_19 (out, din, enable, reset_l, clk) ;
    output  [18:0]  out;
    input   [18:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);

endmodule 


module ff_sre_20 (out, din, enable, reset_l, clk) ;
    output  [19:0]  out;
    input   [19:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);

endmodule 


module ff_sre_21 (out, din, enable, reset_l, clk) ;
    output  [20:0]  out;
    input   [20:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);

endmodule 


module ff_sre_22 (out, din, enable, reset_l, clk) ;
    output  [21:0]  out;
    input   [21:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);

endmodule 


module ff_sre_23 (out, din, enable, reset_l, clk) ;
    output  [22:0]  out;
    input   [22:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);

endmodule 


module ff_sre_24 (out, din, enable, reset_l, clk) ;
    output  [23:0]  out;
    input   [23:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);

endmodule 


module ff_sre_25 (out, din, enable, reset_l, clk) ;
    output  [24:0]  out;
    input   [24:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);

endmodule 


module ff_sre_26 (out, din, enable, reset_l, clk) ;
    output  [25:0]  out;
    input   [25:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);

endmodule 


module ff_sre_27 (out, din, enable, reset_l, clk) ;
    output  [26:0]  out;
    input   [26:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);

endmodule 


module ff_sre_28 (out, din, enable, reset_l, clk) ;
    output  [27:0]  out;
    input   [27:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);
    ff_sre    ff_sre_27(out[27], din[27], enable, reset_l, clk);

endmodule 


module ff_sre_29 (out, din, enable, reset_l, clk) ;
    output  [28:0]  out;
    input   [28:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);
    ff_sre    ff_sre_27(out[27], din[27], enable, reset_l, clk);
    ff_sre    ff_sre_28(out[28], din[28], enable, reset_l, clk);

endmodule 


module ff_sre_30 (out, din, enable, reset_l, clk) ;
    output  [29:0]  out;
    input   [29:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);
    ff_sre    ff_sre_27(out[27], din[27], enable, reset_l, clk);
    ff_sre    ff_sre_28(out[28], din[28], enable, reset_l, clk);
    ff_sre    ff_sre_29(out[29], din[29], enable, reset_l, clk);

endmodule 


module ff_sre_31 (out, din, enable, reset_l, clk) ;
    output  [30:0]  out;
    input   [30:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);
    ff_sre    ff_sre_27(out[27], din[27], enable, reset_l, clk);
    ff_sre    ff_sre_28(out[28], din[28], enable, reset_l, clk);
    ff_sre    ff_sre_29(out[29], din[29], enable, reset_l, clk);
    ff_sre    ff_sre_30(out[30], din[30], enable, reset_l, clk);

endmodule 


module ff_sre_32 (out, din, enable, reset_l, clk) ;
    output  [31:0]  out;
    input   [31:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);
    ff_sre    ff_sre_27(out[27], din[27], enable, reset_l, clk);
    ff_sre    ff_sre_28(out[28], din[28], enable, reset_l, clk);
    ff_sre    ff_sre_29(out[29], din[29], enable, reset_l, clk);
    ff_sre    ff_sre_30(out[30], din[30], enable, reset_l, clk);
    ff_sre    ff_sre_31(out[31], din[31], enable, reset_l, clk);

endmodule 


module ff_sre_40 (out, din, enable, reset_l, clk) ;
    output  [39:0]  out;
    input   [39:0]  din;
    input           clk;
    input           reset_l;
    input           enable;

    ff_sre    ff_sre_0(out[0], din[0], enable, reset_l, clk);
    ff_sre    ff_sre_1(out[1], din[1], enable, reset_l, clk);
    ff_sre    ff_sre_2(out[2], din[2], enable, reset_l, clk);
    ff_sre    ff_sre_3(out[3], din[3], enable, reset_l, clk);
    ff_sre    ff_sre_4(out[4], din[4], enable, reset_l, clk);
    ff_sre    ff_sre_5(out[5], din[5], enable, reset_l, clk);
    ff_sre    ff_sre_6(out[6], din[6], enable, reset_l, clk);
    ff_sre    ff_sre_7(out[7], din[7], enable, reset_l, clk);
    ff_sre    ff_sre_8(out[8], din[8], enable, reset_l, clk);
    ff_sre    ff_sre_9(out[9], din[9], enable, reset_l, clk);
    ff_sre    ff_sre_10(out[10], din[10], enable, reset_l, clk);
    ff_sre    ff_sre_11(out[11], din[11], enable, reset_l, clk);
    ff_sre    ff_sre_12(out[12], din[12], enable, reset_l, clk);
    ff_sre    ff_sre_13(out[13], din[13], enable, reset_l, clk);
    ff_sre    ff_sre_14(out[14], din[14], enable, reset_l, clk);
    ff_sre    ff_sre_15(out[15], din[15], enable, reset_l, clk);
    ff_sre    ff_sre_16(out[16], din[16], enable, reset_l, clk);
    ff_sre    ff_sre_17(out[17], din[17], enable, reset_l, clk);
    ff_sre    ff_sre_18(out[18], din[18], enable, reset_l, clk);
    ff_sre    ff_sre_19(out[19], din[19], enable, reset_l, clk);
    ff_sre    ff_sre_20(out[20], din[20], enable, reset_l, clk);
    ff_sre    ff_sre_21(out[21], din[21], enable, reset_l, clk);
    ff_sre    ff_sre_22(out[22], din[22], enable, reset_l, clk);
    ff_sre    ff_sre_23(out[23], din[23], enable, reset_l, clk);
    ff_sre    ff_sre_24(out[24], din[24], enable, reset_l, clk);
    ff_sre    ff_sre_25(out[25], din[25], enable, reset_l, clk);
    ff_sre    ff_sre_26(out[26], din[26], enable, reset_l, clk);
    ff_sre    ff_sre_27(out[27], din[27], enable, reset_l, clk);
    ff_sre    ff_sre_28(out[28], din[28], enable, reset_l, clk);
    ff_sre    ff_sre_29(out[29], din[29], enable, reset_l, clk);
    ff_sre    ff_sre_30(out[30], din[30], enable, reset_l, clk);
    ff_sre    ff_sre_31(out[31], din[31], enable, reset_l, clk);
    ff_sre    ff_sre_32(out[32], din[32], enable, reset_l, clk);
    ff_sre    ff_sre_33(out[33], din[33], enable, reset_l, clk);
    ff_sre    ff_sre_34(out[34], din[34], enable, reset_l, clk);
    ff_sre    ff_sre_35(out[35], din[35], enable, reset_l, clk);
    ff_sre    ff_sre_36(out[36], din[36], enable, reset_l, clk);
    ff_sre    ff_sre_37(out[37], din[37], enable, reset_l, clk);
    ff_sre    ff_sre_38(out[38], din[38], enable, reset_l, clk);
    ff_sre    ff_sre_39(out[39], din[39], enable, reset_l, clk);

endmodule


module mj_s_ff_snre_d_33 (out, din, lenable, reset_l,clk);
    output  [32:0]  out;
    input   [32:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_23(.out(out[23]), .in(din[23]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_24(.out(out[24]), .in(din[24]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_25(.out(out[25]), .in(din[25]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_26(.out(out[26]), .in(din[26]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_27(.out(out[27]), .in(din[27]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_28(.out(out[28]), .in(din[28]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_29(.out(out[29]), .in(din[29]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_30(.out(out[30]), .in(din[30]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_31(.out(out[31]), .in(din[31]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_32(.out(out[32]), .in(din[32]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snre_d_38 (out, din, lenable, reset_l,clk);
    output  [37:0]  out;
    input   [37:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_23(.out(out[23]), .in(din[23]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_24(.out(out[24]), .in(din[24]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_25(.out(out[25]), .in(din[25]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_26(.out(out[26]), .in(din[26]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_27(.out(out[27]), .in(din[27]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_28(.out(out[28]), .in(din[28]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_29(.out(out[29]), .in(din[29]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_30(.out(out[30]), .in(din[30]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_31(.out(out[31]), .in(din[31]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_32(.out(out[32]), .in(din[32]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_33(.out(out[33]), .in(din[33]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_34(.out(out[34]), .in(din[34]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_35(.out(out[35]), .in(din[35]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_36(.out(out[36]), .in(din[36]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_37(.out(out[37]), .in(din[37]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 

module mj_s_ff_snre_d_64 (out, din, lenable, reset_l,clk);
    output  [63:0]  out;
    input   [63:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_23(.out(out[23]), .in(din[23]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_24(.out(out[24]), .in(din[24]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_25(.out(out[25]), .in(din[25]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_26(.out(out[26]), .in(din[26]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_27(.out(out[27]), .in(din[27]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_28(.out(out[28]), .in(din[28]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_29(.out(out[29]), .in(din[29]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_30(.out(out[30]), .in(din[30]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_31(.out(out[31]), .in(din[31]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_32(.out(out[32]), .in(din[32]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_33(.out(out[33]), .in(din[33]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_34(.out(out[34]), .in(din[34]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_35(.out(out[35]), .in(din[35]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_36(.out(out[36]), .in(din[36]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_37(.out(out[37]), .in(din[37]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_38(.out(out[38]), .in(din[38]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_39(.out(out[39]), .in(din[39]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_40(.out(out[40]), .in(din[40]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_41(.out(out[41]), .in(din[41]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_42(.out(out[42]), .in(din[42]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_43(.out(out[43]), .in(din[43]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_44(.out(out[44]), .in(din[44]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_45(.out(out[45]), .in(din[45]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_46(.out(out[46]), .in(din[46]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_47(.out(out[47]), .in(din[47]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_48(.out(out[48]), .in(din[48]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_49(.out(out[49]), .in(din[49]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_50(.out(out[50]), .in(din[50]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_51(.out(out[51]), .in(din[51]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_52(.out(out[52]), .in(din[52]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_53(.out(out[53]), .in(din[53]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_54(.out(out[54]), .in(din[54]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_55(.out(out[55]), .in(din[55]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_56(.out(out[56]), .in(din[56]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_57(.out(out[57]), .in(din[57]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_58(.out(out[58]), .in(din[58]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_59(.out(out[59]), .in(din[59]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_60(.out(out[60]), .in(din[60]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_61(.out(out[61]), .in(din[61]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_62(.out(out[62]), .in(din[62]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_63(.out(out[63]), .in(din[63]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_2 (out, din, lenable, reset_l,clk);
    output  [1:0]  out;
    input   [1:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;
 
    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
 
endmodule


module mj_s_ff_snre_d_3 (out, din, lenable, reset_l,clk);
    output  [2:0]  out;
    input   [2:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;
 
    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
 
endmodule

module mj_s_ff_snre_d_4 (out, din, lenable, reset_l,clk);
    output  [3:0]  out;
    input   [3:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;
 
    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule


module mj_s_ff_snre_d_18 (out, din, lenable, reset_l,clk);
    output  [17:0]  out;
    input   [17:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 


module mj_s_ff_snre_d_28 (out, din, lenable, reset_l,clk);
    output  [27:0]  out;
    input   [27:0]  din;
    input           lenable;
    input           clk;
    input           reset_l;

    mj_s_ff_snre_d    mj_s_ff_snre_d_0(.out(out[0]), .in(din[0]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_1(.out(out[1]), .in(din[1]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_2(.out(out[2]), .in(din[2]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_3(.out(out[3]), .in(din[3]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_4(.out(out[4]), .in(din[4]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_5(.out(out[5]), .in(din[5]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_6(.out(out[6]), .in(din[6]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_7(.out(out[7]), .in(din[7]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_8(.out(out[8]), .in(din[8]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_9(.out(out[9]), .in(din[9]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_10(.out(out[10]), .in(din[10]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_11(.out(out[11]), .in(din[11]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_12(.out(out[12]), .in(din[12]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_13(.out(out[13]), .in(din[13]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_14(.out(out[14]), .in(din[14]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_15(.out(out[15]), .in(din[15]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_16(.out(out[16]), .in(din[16]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_17(.out(out[17]), .in(din[17]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_18(.out(out[18]), .in(din[18]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_19(.out(out[19]), .in(din[19]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_20(.out(out[20]), .in(din[20]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_21(.out(out[21]), .in(din[21]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_22(.out(out[22]), .in(din[22]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_23(.out(out[23]), .in(din[23]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_24(.out(out[24]), .in(din[24]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_25(.out(out[25]), .in(din[25]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_26(.out(out[26]), .in(din[26]), .lenable(lenable), .reset_l(reset_l),.clk(clk));
    mj_s_ff_snre_d    mj_s_ff_snre_d_27(.out(out[27]), .in(din[27]), .lenable(lenable), .reset_l(reset_l),.clk(clk));

endmodule 

module ff_s_33 (out, din, clk) ;
output [32:0]  out;
input  [32:0]  din;
input          clk;
 
    ff_s    ff_s_0(out[0], din[0], clk);
    ff_s    ff_s_1(out[1], din[1], clk);
    ff_s    ff_s_2(out[2], din[2], clk);
    ff_s    ff_s_3(out[3], din[3], clk);
    ff_s    ff_s_4(out[4], din[4], clk);
    ff_s    ff_s_5(out[5], din[5], clk);
    ff_s    ff_s_6(out[6], din[6], clk);
    ff_s    ff_s_7(out[7], din[7], clk);
    ff_s    ff_s_8(out[8], din[8], clk);
    ff_s    ff_s_9(out[9], din[9], clk);
    ff_s    ff_s_10(out[10], din[10], clk);
    ff_s    ff_s_11(out[11], din[11], clk);
    ff_s    ff_s_12(out[12], din[12], clk);
    ff_s    ff_s_13(out[13], din[13], clk);
    ff_s    ff_s_14(out[14], din[14], clk);
    ff_s    ff_s_15(out[15], din[15], clk);
    ff_s    ff_s_16(out[16], din[16], clk);
    ff_s    ff_s_17(out[17], din[17], clk);
    ff_s    ff_s_18(out[18], din[18], clk);
    ff_s    ff_s_19(out[19], din[19], clk);
    ff_s    ff_s_20(out[20], din[20], clk);
    ff_s    ff_s_21(out[21], din[21], clk);
    ff_s    ff_s_22(out[22], din[22], clk);
    ff_s    ff_s_23(out[23], din[23], clk);
    ff_s    ff_s_24(out[24], din[24], clk);
    ff_s    ff_s_25(out[25], din[25], clk);
    ff_s    ff_s_26(out[26], din[26], clk);
    ff_s    ff_s_27(out[27], din[27], clk);
    ff_s    ff_s_28(out[28], din[28], clk);
    ff_s    ff_s_29(out[29], din[29], clk);
    ff_s    ff_s_30(out[30], din[30], clk);
    ff_s    ff_s_31(out[31], din[31], clk);
    ff_s    ff_s_32(out[32], din[32], clk);
 
endmodule


module ff_drv ( in,out );
input in;
output out;

assign out = in;

endmodule

module ff_drva ( in,out );
input in;
output out;

assign out = in;

endmodule
