/****************************************************************
 ---------------------------------------------------------------
     Copyright 1999 Sun Microsystems, Inc., 901 San Antonio
     Road, Palo Alto, CA 94303, U.S.A.  All Rights Reserved.
     The contents of this file are subject to the current
     version of the Sun Community Source License, picoJava-II
     Core ("the License").  You may not use this file except
     in compliance with the License.  You may obtain a copy
     of the License by searching for "Sun Community Source
     License" on the World Wide Web at http://www.sun.com.
     See the License for the rights, obligations, and
     limitations governing use of the contents of this file.

     Sun, Sun Microsystems, the Sun logo, and all Sun-based
     trademarks and logos, Java, picoJava, and all Java-based
     trademarks and logos are trademarks or registered trademarks 
     of Sun Microsystems, Inc. in the United States and other
     countries.
 ----------------------------------------------------------------
******************************************************************/
                                                  
module ieu_rom (nxt_ucode_cnt,rom_data);          
                                                  
input    [8:0] nxt_ucode_cnt;                     
output  [79:0] rom_data;
                                                  
reg     [79:0] rom_data;
                                                  
/********* Megacell Format **********             
reg     [79:0] mem [511:0];
                                                  
// synopsys translate_off                         
                                                  
initial $readmemh(                                
"picoJava-II/design/iu/ucode/rtl/ieu_rom.data",mem);	// This path needs to be modified based on it's 
						// location.
                                                  
  always @(nxt_ucode_cnt) begin                   
    rom_data = mem[nxt_ucode_cnt];                
  end                                             
                                                  
// synopsys translate_on                          
********** Megacell Format *********/             
                                                  
                                                  
/********* Case    Format **********/             
  always @(nxt_ucode_cnt) begin                   
    case (nxt_ucode_cnt)                          
      9'd000:  rom_data =  80'h00000400000000000000;
      9'd001:  rom_data =  80'h01e2045ca0002780555d;
      9'd002:  rom_data =  80'h00000400000000000000;
      9'd003:  rom_data =  80'h00e204000000000020b8;
      9'd004:  rom_data =  80'h03020442c02666085759;
      9'd005:  rom_data =  80'h00000400000000020000;
      9'd006:  rom_data =  80'h000204000002200002b8;
      9'd007:  rom_data =  80'h00000401203226020959;
      9'd008:  rom_data =  80'h00c604013c0002012b39;
      9'd009:  rom_data =  80'h03020442c02666085759;
      9'd010:  rom_data =  80'h00000400000000020000;
      9'd011:  rom_data =  80'h000204000002200002b8;
      9'd012:  rom_data =  80'h00000419203226020959;
      9'd013:  rom_data =  80'h00c604013c0002012b19;
      9'd014:  rom_data =  80'h03020442c02666085759;
      9'd015:  rom_data =  80'h00000400000000020000;
      9'd016:  rom_data =  80'h000204000002200002b8;
      9'd017:  rom_data =  80'h00000421203226020959;
      9'd018:  rom_data =  80'h00c204013c0002012ab9;
      9'd019:  rom_data =  80'h03020442c02666085759;
      9'd020:  rom_data =  80'h00000400000000020000;
      9'd021:  rom_data =  80'h000204000002200002b8;
      9'd022:  rom_data =  80'h00000429203226020979;
      9'd023:  rom_data =  80'h00c204013c0002010ab9;
      9'd024:  rom_data =  80'h00c2045c000006002b55;
      9'd025:  rom_data =  80'h0000043401bc66000001;
      9'd026:  rom_data =  80'h00080400014000000000;
      9'd027:  rom_data =  80'h01020465a00026085559;
      9'd028:  rom_data =  80'h00000400000000000000;
      9'd029:  rom_data =  80'h000204591800260202b9;
      9'd030:  rom_data =  80'h00000401422026000ad9;
      9'd031:  rom_data =  80'h000404013c000a0326b9;
      9'd032:  rom_data =  80'h0000043401bc66000001;
      9'd033:  rom_data =  80'h00080400014000000000;
      9'd034:  rom_data =  80'h01020465a00026085559;
      9'd035:  rom_data =  80'h00000400000000000000;
      9'd036:  rom_data =  80'h000204591800260202b9;
      9'd037:  rom_data =  80'h00000419422026000ad9;
      9'd038:  rom_data =  80'h000404013c000a0326b9;
      9'd039:  rom_data =  80'h0000043401bc66000001;
      9'd040:  rom_data =  80'h00080400014000000000;
      9'd041:  rom_data =  80'h01020465a00026085559;
      9'd042:  rom_data =  80'h00000400000000000000;
      9'd043:  rom_data =  80'h000204591800260202b9;
      9'd044:  rom_data =  80'h00000421422026000ad9;
      9'd045:  rom_data =  80'h000404013c000a0326b9;
      9'd046:  rom_data =  80'h00000434000ca6000001;
      9'd047:  rom_data =  80'h00080459014022000001;
      9'd048:  rom_data =  80'h010a0465a00026085559;
      9'd049:  rom_data =  80'h00000400000440000000;
      9'd050:  rom_data =  80'h000204591800260202b9;
      9'd051:  rom_data =  80'h000004010224660012db;
      9'd052:  rom_data =  80'h000404013c000a0306b9;
      9'd053:  rom_data =  80'h00040400000010002758;
      9'd054:  rom_data =  80'h00022000000000000c78;
      9'd055:  rom_data =  80'h000004340210860009d1;
      9'd056:  rom_data =  80'h0002040000c220000158;
      9'd057:  rom_data =  80'h00020453003006000759;
      9'd058:  rom_data =  80'h00000401161044000811;
      9'd059:  rom_data =  80'h00020680800120000750;
      9'd060:  rom_data =  80'h00a00409e82226000751;
      9'd061:  rom_data =  80'h004204d9e0002a000bf9;
      9'd062:  rom_data =  80'h006005d9000022000001;
      9'd063:  rom_data =  80'h00800559200022000001;
      9'd064:  rom_data =  80'h00a00600e00008002000;
      9'd065:  rom_data =  80'h00022000000000000c78;
      9'd066:  rom_data =  80'h000004340210860009d1;
      9'd067:  rom_data =  80'h0002040000c220000178;
      9'd068:  rom_data =  80'h00020453003006000751;
      9'd069:  rom_data =  80'h00020409e82026000771;
      9'd070:  rom_data =  80'h00080401161044000811;
      9'd071:  rom_data =  80'h01000400000000004000;
      9'd072:  rom_data =  80'h00000680800120000000;
      9'd073:  rom_data =  80'h00a00400000220000750;
      9'd074:  rom_data =  80'h004204d9e0002a000bf9;
      9'd075:  rom_data =  80'h006005d9000022000001;
      9'd076:  rom_data =  80'h00800559200022000001;
      9'd077:  rom_data =  80'h00a00600e00008002000;
      9'd078:  rom_data =  80'h00000400022220000838;
      9'd079:  rom_data =  80'h00080400000000000000;
      9'd080:  rom_data =  80'h010204000000000054b8;
      9'd081:  rom_data =  80'h000004000210000009d0;
      9'd082:  rom_data =  80'h00020400000000000458;
      9'd083:  rom_data =  80'h00000453003006000001;
      9'd084:  rom_data =  80'h0002040000c220000158;
      9'd085:  rom_data =  80'h00020400000000000750;
      9'd086:  rom_data =  80'h00000401161044000811;
      9'd087:  rom_data =  80'h00000680800120000000;
      9'd088:  rom_data =  80'h00a00400000220000750;
      9'd089:  rom_data =  80'h004204d9e0002a000bf9;
      9'd090:  rom_data =  80'h006005d9000022000001;
      9'd091:  rom_data =  80'h00800559200022000001;
      9'd092:  rom_data =  80'h00a00600e00008002000;
      9'd093:  rom_data =  80'h00022000000000000c78;
      9'd094:  rom_data =  80'h000004000210000009d0;
      9'd095:  rom_data =  80'h00020400000000000178;
      9'd096:  rom_data =  80'h00000400000000000000;
      9'd097:  rom_data =  80'h0000040ce02026000001;
      9'd098:  rom_data =  80'h00080417e03006000001;
      9'd099:  rom_data =  80'h010204000000000054b8;
      9'd100:  rom_data =  80'h00000427403006000001;
      9'd101:  rom_data =  80'h00020400000000000498;
      9'd102:  rom_data =  80'h00000453003006000001;
      9'd103:  rom_data =  80'h0002040000c220000158;
      9'd104:  rom_data =  80'h00020400000000000750;
      9'd105:  rom_data =  80'h00000401161044000811;
      9'd106:  rom_data =  80'h00000680800120000000;
      9'd107:  rom_data =  80'h00a00400000220000750;
      9'd108:  rom_data =  80'h004204d9e0002a000bf9;
      9'd109:  rom_data =  80'h006005d9000022000001;
      9'd110:  rom_data =  80'h00800559200022000001;
      9'd111:  rom_data =  80'h00a00600e00008002000;
      9'd112:  rom_data =  80'h00001073000022000001;
      9'd113:  rom_data =  80'h0008047f003046000001;
      9'd114:  rom_data =  80'h00020400000000001298;
      9'd115:  rom_data =  80'h00000459043006000001;
      9'd116:  rom_data =  80'h00020400000000000098;
      9'd117:  rom_data =  80'h0000047f003006000001;
      9'd118:  rom_data =  80'h000204000000000001f8;
      9'd119:  rom_data =  80'h00000400023000000a78;
      9'd120:  rom_data =  80'h00020400000000000298;
      9'd121:  rom_data =  80'h000004340210860009d1;
      9'd122:  rom_data =  80'h0002040000c220000178;
      9'd123:  rom_data =  80'h00020453003006000751;
      9'd124:  rom_data =  80'h00020409e82026000771;
      9'd125:  rom_data =  80'h00080401161044000811;
      9'd126:  rom_data =  80'h01000400000000004000;
      9'd127:  rom_data =  80'h00000680800120000000;
      9'd128:  rom_data =  80'h00a00400000220000750;
      9'd129:  rom_data =  80'h004204d9e0002a000bf9;
      9'd130:  rom_data =  80'h006005d9000022000001;
      9'd131:  rom_data =  80'h00800559200022000001;
      9'd132:  rom_data =  80'h00a00600e00008002000;
      9'd133:  rom_data =  80'h00001073002002000001;
      9'd134:  rom_data =  80'h00001280200220000cb8;
      9'd135:  rom_data =  80'h00080400000220000770;
      9'd136:  rom_data =  80'h00080480a00220000758;
      9'd137:  rom_data =  80'h00080580a00220000770;
      9'd138:  rom_data =  80'h00080700012000000000;
      9'd139:  rom_data =  80'h00000500200000000000;
      9'd140:  rom_data =  80'h00000600a00000002000;
      9'd141:  rom_data =  80'h00001073002002000001;
      9'd142:  rom_data =  80'h00001280213220000cb8;
      9'd143:  rom_data =  80'h00080400000220000770;
      9'd144:  rom_data =  80'h00080480a00220000758;
      9'd145:  rom_data =  80'h000809dba00262000771;
      9'd146:  rom_data =  80'h000806d9852026000001;
      9'd147:  rom_data =  80'h00a00500200000000000;
      9'd148:  rom_data =  80'h00000600a00000002000;
      9'd149:  rom_data =  80'h00001073002002000001;
      9'd150:  rom_data =  80'h00001280213220000cb8;
      9'd151:  rom_data =  80'h0008040001c220000770;
      9'd152:  rom_data =  80'h00080480a00220000758;
      9'd153:  rom_data =  80'h000809e3a00262000771;
      9'd154:  rom_data =  80'h000806d9852026000001;
      9'd155:  rom_data =  80'h00a00559200026000001;
      9'd156:  rom_data =  80'h00a00600a00008002000;
      9'd157:  rom_data =  80'h00000484c23046000d1a;
      9'd158:  rom_data =  80'h00400564800006000005;
      9'd159:  rom_data =  80'h00a0045c000006002005;
      9'd160:  rom_data =  80'h00000480a00000000000;
      9'd161:  rom_data =  80'h00000700000000000000;
      9'd162:  rom_data =  80'h00000500c00000000000;
      9'd163:  rom_data =  80'h00000400000000002000;
      9'd164:  rom_data =  80'h000008ecc22026000d51;
      9'd165:  rom_data =  80'h00080ab3213026000001;
      9'd166:  rom_data =  80'h00a00500a00000000000;
      9'd167:  rom_data =  80'h00000400000000002000;
      9'd168:  rom_data =  80'h0000086c022026000d71;
      9'd169:  rom_data =  80'h000806d9213026000001;
      9'd170:  rom_data =  80'h000808dba00022000001;
      9'd171:  rom_data =  80'h00a00559a1b026000001;
      9'd172:  rom_data =  80'h00a00400000000002000;
      9'd173:  rom_data =  80'h0000045e022026000cb9;
      9'd174:  rom_data =  80'h000204000000000006b8;
      9'd175:  rom_data =  80'h00020400000220000758;
      9'd176:  rom_data =  80'h00020401341226000759;
      9'd177:  rom_data =  80'h00000402e03a62000759;
      9'd178:  rom_data =  80'h00000480023000000a98;
      9'd179:  rom_data =  80'h00000402900222200699;
      9'd180:  rom_data =  80'h00000402f00224300699;
      9'd181:  rom_data =  80'h000204000000000006b8;
      9'd182:  rom_data =  80'h00000400000000000000;
      9'd183:  rom_data =  80'h00000401342006000001;
      9'd184:  rom_data =  80'h00000480200000002000;
      9'd185:  rom_data =  80'h010204000000001014b8;
      9'd186:  rom_data =  80'h00022000000000000c78;
      9'd187:  rom_data =  80'h00020400000000000570;
      9'd188:  rom_data =  80'h00000400009000000000;
      9'd189:  rom_data =  80'h00000401140044000001;
      9'd190:  rom_data =  80'h0200040080000000a000;
      9'd191:  rom_data =  80'h010204000000001014b8;
      9'd192:  rom_data =  80'h00022000000000000c78;
      9'd193:  rom_data =  80'h00020447003006000571;
      9'd194:  rom_data =  80'h00000400009000000000;
      9'd195:  rom_data =  80'h00000401140044000001;
      9'd196:  rom_data =  80'h0200045c800026008001;
      9'd197:  rom_data =  80'h00a00400000000002000;
      9'd198:  rom_data =  80'h00001000000220000dd0;
      9'd199:  rom_data =  80'h00080400000000000000;
      9'd200:  rom_data =  80'h00000480a00000002000;
      9'd201:  rom_data =  80'h00001073000022000001;
      9'd202:  rom_data =  80'h0008047f003226000959;
      9'd203:  rom_data =  80'h00c20400000000003298;
      9'd204:  rom_data =  80'h00a0045c000c9e000005;
      9'd205:  rom_data =  80'h00a0046400023600099d;
      9'd206:  rom_data =  80'h00a00400000018002000;
      9'd207:  rom_data =  80'h00a0045c021c9e0009bd;
      9'd208:  rom_data =  80'h00b0046401423600099d;
      9'd209:  rom_data =  80'h00a00400000138000000;
      9'd210:  rom_data =  80'h00a00400000008002000;
      9'd211:  rom_data =  80'h00a0045c000c9e000005;
      9'd212:  rom_data =  80'h00a00464000016002005;
      9'd213:  rom_data =  80'h00a0045c021c9e0009dd;
      9'd214:  rom_data =  80'h00b00464014016000005;
      9'd215:  rom_data =  80'h00a0046c00023e0009bd;
      9'd216:  rom_data =  80'h00a00400000128000000;
      9'd217:  rom_data =  80'h00a00400000010002000;
      9'd218:  rom_data =  80'h00a0045c021ebe0009dd;
      9'd219:  rom_data =  80'h00b00464014016000005;
      9'd220:  rom_data =  80'h00a0046c02101e00075d;
      9'd221:  rom_data =  80'h00b004000002280009b8;
      9'd222:  rom_data =  80'h00a00400000138000000;
      9'd223:  rom_data =  80'h00a00400000010002000;
      9'd224:  rom_data =  80'h00a00464000c9e000005;
      9'd225:  rom_data =  80'h00a0045c000036002005;
      9'd226:  rom_data =  80'h00c2205c023006002c5d;
      9'd227:  rom_data =  80'h00c2205c023006002c7d;
      9'd228:  rom_data =  80'h00c2205c023006000c7d;
      9'd229:  rom_data =  80'h00c20464000006002b5d;
      9'd230:  rom_data =  80'h01c2045ca2100700547d;
      9'd231:  rom_data =  80'h00020400000220001558;
      9'd232:  rom_data =  80'h00000401000024000001;
      9'd233:  rom_data =  80'h00c2045c00000600261d;
      9'd234:  rom_data =  80'h03040400c21019005678;
      9'd235:  rom_data =  80'h00020400000220001758;
      9'd236:  rom_data =  80'h00000401000024000001;
      9'd237:  rom_data =  80'h00040400000018002618;
      9'd238:  rom_data =  80'h01c2045ca2122684547d;
      9'd239:  rom_data =  80'h00c2046400002600275d;
      9'd240:  rom_data =  80'h00020400000220001558;
      9'd241:  rom_data =  80'h00000401000024000001;
      9'd242:  rom_data =  80'h00c2045c00022600061d;
      9'd243:  rom_data =  80'h00c2046400000600275d;
      9'd244:  rom_data =  80'h0304045cc2103a8c5679;
      9'd245:  rom_data =  80'h00080400000120000000;
      9'd246:  rom_data =  80'h00040400000018002758;
      9'd247:  rom_data =  80'h000a0400014220001758;
      9'd248:  rom_data =  80'h00000401000024000001;
      9'd249:  rom_data =  80'h00040400000228000618;
      9'd250:  rom_data =  80'h00040400000018002758;
      9'd251:  rom_data =  80'h00022000000000000c78;
      9'd252:  rom_data =  80'h0000045c000026000001;
      9'd253:  rom_data =  80'h00c204000000000022b8;
      9'd254:  rom_data =  80'h00022000000000000c78;
      9'd255:  rom_data =  80'h00000400000000000000;
      9'd256:  rom_data =  80'h000404000000180022b8;
      9'd257:  rom_data =  80'h00022000000000000c78;
      9'd258:  rom_data =  80'h0000045c000026000001;
      9'd259:  rom_data =  80'h00c204640230260002b9;
      9'd260:  rom_data =  80'h00c20400000000002b58;
      9'd261:  rom_data =  80'h00022000000c80000c78;
      9'd262:  rom_data =  80'h00000400000000000000;
      9'd263:  rom_data =  80'h000404000000180002b8;
      9'd264:  rom_data =  80'h00040400000010002358;
      9'd265:  rom_data =  80'h03048000d21019405678;
      9'd266:  rom_data =  80'h00020400000220001758;
      9'd267:  rom_data =  80'h00000401000024000001;
      9'd268:  rom_data =  80'h00040400000018002618;
      9'd269:  rom_data =  80'h00022000000c80000c78;
      9'd270:  rom_data =  80'h00000400000000000000;
      9'd271:  rom_data =  80'h00048000f000184022b8;
      9'd272:  rom_data =  80'h0000106b002002000001;
      9'd273:  rom_data =  80'h00001280200220000cb8;
      9'd274:  rom_data =  80'h00080400000220000770;
      9'd275:  rom_data =  80'h00080480a00220000758;
      9'd276:  rom_data =  80'h00080580a00220000778;
      9'd277:  rom_data =  80'h00080700012000000000;
      9'd278:  rom_data =  80'h00000500200000000000;
      9'd279:  rom_data =  80'h00000780a00000002000;
      9'd280:  rom_data =  80'h00000474023026000cb9;
      9'd281:  rom_data =  80'h00204059024062000eb9;
      9'd282:  rom_data =  80'h00a303e1600022000cb1;
      9'd283:  rom_data =  80'h006005d9800026000001;
      9'd284:  rom_data =  80'h00400480e00000002000;
      9'd285:  rom_data =  80'h0000043401bc66000001;
      9'd286:  rom_data =  80'h00080400014480000000;
      9'd287:  rom_data =  80'h01020465a00026085559;
      9'd288:  rom_data =  80'h00000400000000000000;
      9'd289:  rom_data =  80'h000204591800260202b9;
      9'd290:  rom_data =  80'h00000421422026000ad9;
      9'd291:  rom_data =  80'h000004013c0002030001;
      9'd292:  rom_data =  80'h00048000a800084026b8;
      9'd293:  rom_data =  80'h010204000000001014b8;
      9'd294:  rom_data =  80'h00000400000000000000;
      9'd295:  rom_data =  80'h00000400000000002000;
      9'd296:  rom_data =  80'h00000400000000000000;
      9'd297:  rom_data =  80'h00000400000000000000;
      9'd298:  rom_data =  80'h00000400000000000000;
      9'd299:  rom_data =  80'h00000400000000000000;
      default: rom_data =  80'h00000400000000000000;
    endcase                               
  end // end the always                   
/********* Case    Format **********/     
                                          
endmodule                                 
